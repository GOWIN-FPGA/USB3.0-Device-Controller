module gw_gao(
    \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/in_data[31] ,
    \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/in_data[30] ,
    \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/in_data[29] ,
    \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/in_data[28] ,
    \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/in_data[27] ,
    \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/in_data[26] ,
    \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/in_data[25] ,
    \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/in_data[24] ,
    \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/in_data[23] ,
    \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/in_data[22] ,
    \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/in_data[21] ,
    \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/in_data[20] ,
    \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/in_data[19] ,
    \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/in_data[18] ,
    \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/in_data[17] ,
    \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/in_data[16] ,
    \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/in_data[15] ,
    \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/in_data[14] ,
    \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/in_data[13] ,
    \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/in_data[12] ,
    \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/in_data[11] ,
    \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/in_data[10] ,
    \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/in_data[9] ,
    \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/in_data[8] ,
    \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/in_data[7] ,
    \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/in_data[6] ,
    \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/in_data[5] ,
    \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/in_data[4] ,
    \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/in_data[3] ,
    \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/in_data[2] ,
    \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/in_data[1] ,
    \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/in_data[0] ,
    \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/in_datak[3] ,
    \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/in_datak[2] ,
    \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/in_datak[1] ,
    \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/in_datak[0] ,
    \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/in_active ,
    \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/outp_data[31] ,
    \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/outp_data[30] ,
    \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/outp_data[29] ,
    \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/outp_data[28] ,
    \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/outp_data[27] ,
    \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/outp_data[26] ,
    \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/outp_data[25] ,
    \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/outp_data[24] ,
    \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/outp_data[23] ,
    \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/outp_data[22] ,
    \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/outp_data[21] ,
    \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/outp_data[20] ,
    \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/outp_data[19] ,
    \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/outp_data[18] ,
    \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/outp_data[17] ,
    \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/outp_data[16] ,
    \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/outp_data[15] ,
    \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/outp_data[14] ,
    \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/outp_data[13] ,
    \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/outp_data[12] ,
    \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/outp_data[11] ,
    \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/outp_data[10] ,
    \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/outp_data[9] ,
    \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/outp_data[8] ,
    \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/outp_data[7] ,
    \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/outp_data[6] ,
    \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/outp_data[5] ,
    \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/outp_data[4] ,
    \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/outp_data[3] ,
    \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/outp_data[2] ,
    \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/outp_data[1] ,
    \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/outp_data[0] ,
    \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/outp_datak[3] ,
    \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/outp_datak[2] ,
    \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/outp_datak[1] ,
    \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/outp_datak[0] ,
    \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/outp_active ,
    \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/out_stall ,
    \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/enter_u0_cnt[7] ,
    \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/enter_u0_cnt[6] ,
    \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/enter_u0_cnt[5] ,
    \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/enter_u0_cnt[4] ,
    \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/enter_u0_cnt[3] ,
    \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/enter_u0_cnt[2] ,
    \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/enter_u0_cnt[1] ,
    \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/enter_u0_cnt[0] ,
    \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/ltssm_exit_u0 ,
    \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/ltssm_current_state[4] ,
    \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/ltssm_current_state[3] ,
    \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/ltssm_current_state[2] ,
    \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/ltssm_current_state[1] ,
    \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/ltssm_current_state[0] ,
    \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/queue_send_u0_adv ,
    \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/queue_send_u0_portcap ,
    \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/link_cmd_det ,
    \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/send_port_cfg_resp ,
    \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/remote_rx_cred_count[2] ,
    \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/remote_rx_cred_count[1] ,
    \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/remote_rx_cred_count[0] ,
    \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/tx_cred_idx[1] ,
    \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/tx_cred_idx[0] ,
    \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/send_port_cfg_resp_ack ,
    \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/ack_tx_hdr_seq_num[2] ,
    \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/ack_tx_hdr_seq_num[1] ,
    \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/ack_tx_hdr_seq_num[0] ,
    \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/rx_hdr_seq_num[2] ,
    \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/rx_hdr_seq_num[1] ,
    \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/rx_hdr_seq_num[0] ,
    \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/ltssm_enter_u0_by_polling ,
    \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/in_link_command_act ,
    \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/in_link_command_crc_good ,
    \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/in_link_command_latch_act ,
    \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/recv_u0_adv ,
    \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/err_lgood_order ,
    \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/err_lcrd_mismatch ,
    \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/err_lbad_recv ,
    \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/hp_det ,
    \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/in_header_act ,
    \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/hp_crc_good ,
    \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/err_hp_seq ,
    \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/err_lbad ,
    \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/local_rx_cred_count[2] ,
    \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/local_rx_cred_count[1] ,
    \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/local_rx_cred_count[0] ,
    \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/rx_dph ,
    \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/rx_dph_eob ,
    \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/rx_dph_setup ,
    \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/rx_dph_pktpend ,
    \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/rx_dph_endp[3] ,
    \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/rx_dph_endp[2] ,
    \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/rx_dph_endp[1] ,
    \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/rx_dph_endp[0] ,
    \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/rx_dph_seq[4] ,
    \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/rx_dph_seq[3] ,
    \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/rx_dph_seq[2] ,
    \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/rx_dph_seq[1] ,
    \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/rx_dph_seq[0] ,
    \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/rx_dph_len[15] ,
    \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/rx_dph_len[14] ,
    \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/rx_dph_len[13] ,
    \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/rx_dph_len[12] ,
    \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/rx_dph_len[11] ,
    \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/rx_dph_len[10] ,
    \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/rx_dph_len[9] ,
    \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/rx_dph_len[8] ,
    \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/rx_dph_len[7] ,
    \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/rx_dph_len[6] ,
    \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/rx_dph_len[5] ,
    \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/rx_dph_len[4] ,
    \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/rx_dph_len[3] ,
    \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/rx_dph_len[2] ,
    \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/rx_dph_len[1] ,
    \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/rx_dph_len[0] ,
    \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/rx_tp_subtype[3] ,
    \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/rx_tp_subtype[2] ,
    \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/rx_tp_subtype[1] ,
    \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/rx_tp_subtype[0] ,
    \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/rx_tp_endp[3] ,
    \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/rx_tp_endp[2] ,
    \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/rx_tp_endp[1] ,
    \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/rx_tp_endp[0] ,
    \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/rx_tp_nump[4] ,
    \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/rx_tp_nump[3] ,
    \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/rx_tp_nump[2] ,
    \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/rx_tp_nump[1] ,
    \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/rx_tp_nump[0] ,
    \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/rx_tp_seq[4] ,
    \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/rx_tp_seq[3] ,
    \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/rx_tp_seq[2] ,
    \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/rx_tp_seq[1] ,
    \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/rx_tp_seq[0] ,
    \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/rx_tp_stream[15] ,
    \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/rx_tp_stream[14] ,
    \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/rx_tp_stream[13] ,
    \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/rx_tp_stream[12] ,
    \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/rx_tp_stream[11] ,
    \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/rx_tp_stream[10] ,
    \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/rx_tp_stream[9] ,
    \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/rx_tp_stream[8] ,
    \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/rx_tp_stream[7] ,
    \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/rx_tp_stream[6] ,
    \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/rx_tp_stream[5] ,
    \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/rx_tp_stream[4] ,
    \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/rx_tp_stream[3] ,
    \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/rx_tp_stream[2] ,
    \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/rx_tp_stream[1] ,
    \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/rx_tp_stream[0] ,
    \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/rx_tp ,
    \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/rx_tp_retry ,
    \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/rx_tp_pktpend ,
    \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/tx_tp_a_subtype[3] ,
    \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/tx_tp_a_subtype[2] ,
    \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/tx_tp_a_subtype[1] ,
    \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/tx_tp_a_subtype[0] ,
    \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/tx_tp_a_endp[3] ,
    \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/tx_tp_a_endp[2] ,
    \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/tx_tp_a_endp[1] ,
    \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/tx_tp_a_endp[0] ,
    \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/tx_tp_a ,
    \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/tx_tp_a_dir ,
    \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/tx_tp_a_nump[4] ,
    \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/tx_tp_a_nump[3] ,
    \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/tx_tp_a_nump[2] ,
    \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/tx_tp_a_nump[1] ,
    \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/tx_tp_a_nump[0] ,
    \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/tx_tp_a_seq[4] ,
    \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/tx_tp_a_seq[3] ,
    \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/tx_tp_a_seq[2] ,
    \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/tx_tp_a_seq[1] ,
    \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/tx_tp_a_seq[0] ,
    \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/tx_tp_a_stream[15] ,
    \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/tx_tp_a_stream[14] ,
    \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/tx_tp_a_stream[13] ,
    \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/tx_tp_a_stream[12] ,
    \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/tx_tp_a_stream[11] ,
    \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/tx_tp_a_stream[10] ,
    \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/tx_tp_a_stream[9] ,
    \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/tx_tp_a_stream[8] ,
    \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/tx_tp_a_stream[7] ,
    \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/tx_tp_a_stream[6] ,
    \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/tx_tp_a_stream[5] ,
    \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/tx_tp_a_stream[4] ,
    \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/tx_tp_a_stream[3] ,
    \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/tx_tp_a_stream[2] ,
    \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/tx_tp_a_stream[1] ,
    \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/tx_tp_a_stream[0] ,
    \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/tx_tp_a_retry ,
    \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/tx_tp_b_subtype[3] ,
    \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/tx_tp_b_subtype[2] ,
    \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/tx_tp_b_subtype[1] ,
    \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/tx_tp_b_subtype[0] ,
    \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/tx_tp_b_endp[3] ,
    \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/tx_tp_b_endp[2] ,
    \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/tx_tp_b_endp[1] ,
    \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/tx_tp_b_endp[0] ,
    \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/tx_tp_b ,
    \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/tx_tp_b_retry ,
    \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/tx_tp_b_nump[4] ,
    \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/tx_tp_b_nump[3] ,
    \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/tx_tp_b_nump[2] ,
    \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/tx_tp_b_nump[1] ,
    \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/tx_tp_b_nump[0] ,
    \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/tx_tp_c_subtype[3] ,
    \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/tx_tp_c_subtype[2] ,
    \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/tx_tp_c_subtype[1] ,
    \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/tx_tp_c_subtype[0] ,
    \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/tx_tp_c_endp[3] ,
    \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/tx_tp_c_endp[2] ,
    \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/tx_tp_c_endp[1] ,
    \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/tx_tp_c_endp[0] ,
    \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/tx_tp_c ,
    \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/tx_tp_c_retry ,
    \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/tx_tp_c_nump[4] ,
    \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/tx_tp_c_nump[3] ,
    \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/tx_tp_c_nump[2] ,
    \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/tx_tp_c_nump[1] ,
    \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/tx_tp_c_nump[0] ,
    \UserLayer_top_inst/DataTransfer_inst/ep1_in_buf_ready ,
    \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/iu3ep0/req_cnt[7] ,
    \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/iu3ep0/req_cnt[6] ,
    \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/iu3ep0/req_cnt[5] ,
    \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/iu3ep0/req_cnt[4] ,
    \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/iu3ep0/req_cnt[3] ,
    \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/iu3ep0/req_cnt[2] ,
    \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/iu3ep0/req_cnt[1] ,
    \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/iu3ep0/req_cnt[0] ,
    \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/host_requests_data ,
    \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/host_requests_endpt[3] ,
    \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/host_requests_endpt[2] ,
    \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/host_requests_endpt[1] ,
    \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/host_requests_endpt[0] ,
    \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/rx_dpp_start ,
    \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/rx_dpp_done ,
    \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/rx_dpp_crcgood ,
    \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/err_missed_dpp_start ,
    \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/err_missed_dpp_done ,
    \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/tx_dph ,
    \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/tx_dph_eob ,
    \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/tx_dph_dir ,
    \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/tx_dph_endp[3] ,
    \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/tx_dph_endp[2] ,
    \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/tx_dph_endp[1] ,
    \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/tx_dph_endp[0] ,
    \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/tx_dph_seq[4] ,
    \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/tx_dph_seq[3] ,
    \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/tx_dph_seq[2] ,
    \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/tx_dph_seq[1] ,
    \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/tx_dph_seq[0] ,
    \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/tx_dph_len[15] ,
    \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/tx_dph_len[14] ,
    \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/tx_dph_len[13] ,
    \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/tx_dph_len[12] ,
    \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/tx_dph_len[11] ,
    \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/tx_dph_len[10] ,
    \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/tx_dph_len[9] ,
    \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/tx_dph_len[8] ,
    \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/tx_dph_len[7] ,
    \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/tx_dph_len[6] ,
    \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/tx_dph_len[5] ,
    \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/tx_dph_len[4] ,
    \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/tx_dph_len[3] ,
    \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/tx_dph_len[2] ,
    \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/tx_dph_len[1] ,
    \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/tx_dph_len[0] ,
    \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/tx_dpp_ack ,
    \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/tx_dpp_done ,
    \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/ep2_buf_out_nump[4] ,
    \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/ep2_buf_out_nump[3] ,
    \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/ep2_buf_out_nump[2] ,
    \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/ep2_buf_out_nump[1] ,
    \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/ep2_buf_out_nump[0] ,
    \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/burst_in_act ,
    \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/burst_in_stop ,
    \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/do_send_dpp ,
    \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/do_send_dpp_ack ,
    \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/do_send_dpp_eob ,
    \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/crc_hprx_out[15] ,
    \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/crc_hprx_out[14] ,
    \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/crc_hprx_out[13] ,
    \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/crc_hprx_out[12] ,
    \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/crc_hprx_out[11] ,
    \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/crc_hprx_out[10] ,
    \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/crc_hprx_out[9] ,
    \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/crc_hprx_out[8] ,
    \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/crc_hprx_out[7] ,
    \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/crc_hprx_out[6] ,
    \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/crc_hprx_out[5] ,
    \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/crc_hprx_out[4] ,
    \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/crc_hprx_out[3] ,
    \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/crc_hprx_out[2] ,
    \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/crc_hprx_out[1] ,
    \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/crc_hprx_out[0] ,
    \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/crc_hprx_rst ,
    \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/crc_hprx_en ,
    \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/crc_hprx_in[31] ,
    \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/crc_hprx_in[30] ,
    \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/crc_hprx_in[29] ,
    \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/crc_hprx_in[28] ,
    \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/crc_hprx_in[27] ,
    \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/crc_hprx_in[26] ,
    \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/crc_hprx_in[25] ,
    \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/crc_hprx_in[24] ,
    \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/crc_hprx_in[23] ,
    \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/crc_hprx_in[22] ,
    \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/crc_hprx_in[21] ,
    \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/crc_hprx_in[20] ,
    \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/crc_hprx_in[19] ,
    \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/crc_hprx_in[18] ,
    \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/crc_hprx_in[17] ,
    \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/crc_hprx_in[16] ,
    \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/crc_hprx_in[15] ,
    \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/crc_hprx_in[14] ,
    \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/crc_hprx_in[13] ,
    \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/crc_hprx_in[12] ,
    \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/crc_hprx_in[11] ,
    \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/crc_hprx_in[10] ,
    \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/crc_hprx_in[9] ,
    \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/crc_hprx_in[8] ,
    \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/crc_hprx_in[7] ,
    \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/crc_hprx_in[6] ,
    \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/crc_hprx_in[5] ,
    \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/crc_hprx_in[4] ,
    \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/crc_hprx_in[3] ,
    \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/crc_hprx_in[2] ,
    \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/crc_hprx_in[1] ,
    \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/crc_hprx_in[0] ,
    \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/crc_cw3_out[4] ,
    \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/crc_cw3_out[3] ,
    \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/crc_cw3_out[2] ,
    \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/crc_cw3_out[1] ,
    \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/crc_cw3_out[0] ,
    \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/in_header_cw[15] ,
    \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/in_header_cw[14] ,
    \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/in_header_cw[13] ,
    \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/in_header_cw[12] ,
    \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/in_header_cw[11] ,
    \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/in_header_cw[10] ,
    \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/in_header_cw[9] ,
    \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/in_header_cw[8] ,
    \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/in_header_cw[7] ,
    \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/in_header_cw[6] ,
    \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/in_header_cw[5] ,
    \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/in_header_cw[4] ,
    \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/in_header_cw[3] ,
    \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/in_header_cw[2] ,
    \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/in_header_cw[1] ,
    \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/in_header_cw[0] ,
    \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/in_link_command[10] ,
    \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/in_link_command[9] ,
    \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/in_link_command[8] ,
    \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/in_link_command[7] ,
    \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/in_link_command[6] ,
    \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/in_link_command[5] ,
    \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/in_link_command[4] ,
    \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/in_link_command[3] ,
    \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/in_link_command[2] ,
    \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/in_link_command[1] ,
    \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/in_link_command[0] ,
    \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/crc_cw1_out[4] ,
    \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/crc_cw1_out[3] ,
    \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/crc_cw1_out[2] ,
    \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/crc_cw1_out[1] ,
    \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/crc_cw1_out[0] ,
    \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/in_link_command[31] ,
    \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/in_link_command[30] ,
    \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/in_link_command[29] ,
    \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/in_link_command[28] ,
    \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/in_link_command[27] ,
    \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/in_link_command[26] ,
    \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/in_link_command[25] ,
    \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/in_link_command[24] ,
    \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/in_link_command[23] ,
    \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/in_link_command[22] ,
    \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/in_link_command[21] ,
    \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/in_link_command[20] ,
    \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/in_link_command[19] ,
    \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/in_link_command[18] ,
    \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/in_link_command[17] ,
    \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/in_link_command[16] ,
    \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/crc_cw2_out[4] ,
    \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/crc_cw2_out[3] ,
    \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/crc_cw2_out[2] ,
    \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/crc_cw2_out[1] ,
    \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/crc_cw2_out[0] ,
    \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/in_link_command[15] ,
    \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/in_link_command[14] ,
    \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/in_link_command[13] ,
    \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/in_link_command[12] ,
    \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/in_link_command[11] ,
    \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/err_lbad_reg ,
    \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/rx_hdr_seq_num_reg[2] ,
    \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/rx_hdr_seq_num_reg[1] ,
    \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/rx_hdr_seq_num_reg[0] ,
    \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/link_err ,
    \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/tx_lbad_pop ,
    \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/tx_lbad_q[10] ,
    \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/tx_lbad_q[9] ,
    \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/tx_lbad_q[8] ,
    \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/tx_lbad_q[7] ,
    \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/tx_lbad_q[6] ,
    \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/tx_lbad_q[5] ,
    \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/tx_lbad_q[4] ,
    \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/tx_lbad_q[3] ,
    \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/tx_lbad_q[2] ,
    \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/tx_lbad_q[1] ,
    \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/tx_lbad_q[0] ,
    \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/tx_lbad_empty ,
    \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/tx_lbad_act ,
    \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/wait_retry ,
    \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/rx_retry ,
    \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/hp_valid_k_cnt[2] ,
    \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/hp_valid_k_cnt[1] ,
    \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/hp_valid_k_cnt[0] ,
    \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/hp_valid_k[3] ,
    \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/hp_valid_k[2] ,
    \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/hp_valid_k[1] ,
    \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/hp_valid_k[0] ,
    \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/queue_state[2] ,
    \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/queue_state[1] ,
    \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/queue_state[0] ,
    \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/send_dpp_state[3] ,
    \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/send_dpp_state[2] ,
    \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/send_dpp_state[1] ,
    \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/send_dpp_state[0] ,
    \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/tx_link_busy ,
    \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/tx_lcmd_req ,
    \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/tx_hp_req ,
    \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/ltssm_state[4] ,
    \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/ltssm_state[3] ,
    \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/ltssm_state[2] ,
    \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/ltssm_state[1] ,
    \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/ltssm_state[0] ,
    \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/reset_n ,
    \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/ltssm_go_recovery ,
    \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/res_mem_wr_en ,
    \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/res_mem_wr_dat[35] ,
    \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/res_mem_wr_dat[34] ,
    \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/res_mem_wr_dat[33] ,
    \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/res_mem_wr_dat[32] ,
    \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/res_mem_wr_dat[31] ,
    \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/res_mem_wr_dat[30] ,
    \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/res_mem_wr_dat[29] ,
    \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/res_mem_wr_dat[28] ,
    \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/res_mem_wr_dat[27] ,
    \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/res_mem_wr_dat[26] ,
    \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/res_mem_wr_dat[25] ,
    \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/res_mem_wr_dat[24] ,
    \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/res_mem_wr_dat[23] ,
    \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/res_mem_wr_dat[22] ,
    \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/res_mem_wr_dat[21] ,
    \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/res_mem_wr_dat[20] ,
    \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/res_mem_wr_dat[19] ,
    \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/res_mem_wr_dat[18] ,
    \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/res_mem_wr_dat[17] ,
    \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/res_mem_wr_dat[16] ,
    \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/res_mem_wr_dat[15] ,
    \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/res_mem_wr_dat[14] ,
    \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/res_mem_wr_dat[13] ,
    \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/res_mem_wr_dat[12] ,
    \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/res_mem_wr_dat[11] ,
    \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/res_mem_wr_dat[10] ,
    \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/res_mem_wr_dat[9] ,
    \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/res_mem_wr_dat[8] ,
    \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/res_mem_wr_dat[7] ,
    \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/res_mem_wr_dat[6] ,
    \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/res_mem_wr_dat[5] ,
    \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/res_mem_wr_dat[4] ,
    \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/res_mem_wr_dat[3] ,
    \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/res_mem_wr_dat[2] ,
    \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/res_mem_wr_dat[1] ,
    \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/res_mem_wr_dat[0] ,
    \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/res_mem_wr_addr[10] ,
    \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/res_mem_wr_addr[9] ,
    \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/res_mem_wr_addr[8] ,
    \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/res_mem_wr_addr[7] ,
    \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/res_mem_wr_addr[6] ,
    \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/res_mem_wr_addr[5] ,
    \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/res_mem_wr_addr[4] ,
    \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/res_mem_wr_addr[3] ,
    \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/res_mem_wr_addr[2] ,
    \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/res_mem_wr_addr[1] ,
    \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/res_mem_wr_addr[0] ,
    \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/res_mem_wr_pt[1] ,
    \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/res_mem_wr_pt[0] ,
    \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/resend_hp_act ,
    \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/tx_hdr_seq_num_dec[2] ,
    \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/tx_hdr_seq_num_dec[1] ,
    \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/tx_hdr_seq_num_dec[0] ,
    \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/resend_hp_num[4] ,
    \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/resend_hp_num[3] ,
    \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/resend_hp_num[2] ,
    \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/resend_hp_num[1] ,
    \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/resend_hp_num[0] ,
    \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/res_mem_rd_pt[1] ,
    \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/res_mem_rd_pt[0] ,
    \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/res_mem_rd_addr[10] ,
    \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/res_mem_rd_addr[9] ,
    \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/res_mem_rd_addr[8] ,
    \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/res_mem_rd_addr[7] ,
    \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/res_mem_rd_addr[6] ,
    \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/res_mem_rd_addr[5] ,
    \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/res_mem_rd_addr[4] ,
    \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/res_mem_rd_addr[3] ,
    \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/res_mem_rd_addr[2] ,
    \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/res_mem_rd_addr[1] ,
    \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/res_mem_rd_addr[0] ,
    \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/res_mem_rd_en ,
    \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/tx_res_req ,
    \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/tx_res_req_ack ,
    \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/res_mem_rd_dat[35] ,
    \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/res_mem_rd_dat[34] ,
    \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/res_mem_rd_dat[33] ,
    \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/res_mem_rd_dat[32] ,
    \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/res_mem_rd_dat[31] ,
    \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/res_mem_rd_dat[30] ,
    \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/res_mem_rd_dat[29] ,
    \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/res_mem_rd_dat[28] ,
    \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/res_mem_rd_dat[27] ,
    \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/res_mem_rd_dat[26] ,
    \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/res_mem_rd_dat[25] ,
    \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/res_mem_rd_dat[24] ,
    \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/res_mem_rd_dat[23] ,
    \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/res_mem_rd_dat[22] ,
    \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/res_mem_rd_dat[21] ,
    \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/res_mem_rd_dat[20] ,
    \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/res_mem_rd_dat[19] ,
    \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/res_mem_rd_dat[18] ,
    \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/res_mem_rd_dat[17] ,
    \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/res_mem_rd_dat[16] ,
    \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/res_mem_rd_dat[15] ,
    \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/res_mem_rd_dat[14] ,
    \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/res_mem_rd_dat[13] ,
    \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/res_mem_rd_dat[12] ,
    \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/res_mem_rd_dat[11] ,
    \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/res_mem_rd_dat[10] ,
    \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/res_mem_rd_dat[9] ,
    \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/res_mem_rd_dat[8] ,
    \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/res_mem_rd_dat[7] ,
    \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/res_mem_rd_dat[6] ,
    \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/res_mem_rd_dat[5] ,
    \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/res_mem_rd_dat[4] ,
    \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/res_mem_rd_dat[3] ,
    \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/res_mem_rd_dat[2] ,
    \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/res_mem_rd_dat[1] ,
    \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/res_mem_rd_dat[0] ,
    \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/res_mem_rd_dat_val ,
    \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/out_data_5[31] ,
    \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/out_data_5[30] ,
    \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/out_data_5[29] ,
    \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/out_data_5[28] ,
    \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/out_data_5[27] ,
    \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/out_data_5[26] ,
    \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/out_data_5[25] ,
    \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/out_data_5[24] ,
    \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/out_data_5[23] ,
    \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/out_data_5[22] ,
    \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/out_data_5[21] ,
    \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/out_data_5[20] ,
    \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/out_data_5[19] ,
    \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/out_data_5[18] ,
    \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/out_data_5[17] ,
    \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/out_data_5[16] ,
    \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/out_data_5[15] ,
    \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/out_data_5[14] ,
    \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/out_data_5[13] ,
    \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/out_data_5[12] ,
    \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/out_data_5[11] ,
    \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/out_data_5[10] ,
    \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/out_data_5[9] ,
    \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/out_data_5[8] ,
    \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/out_data_5[7] ,
    \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/out_data_5[6] ,
    \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/out_data_5[5] ,
    \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/out_data_5[4] ,
    \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/out_data_5[3] ,
    \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/out_data_5[2] ,
    \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/out_data_5[1] ,
    \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/out_data_5[0] ,
    \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/out_datak_5[3] ,
    \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/out_datak_5[2] ,
    \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/out_datak_5[1] ,
    \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/out_datak_5[0] ,
    \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/out_active_5 ,
    \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/tx_hdr_seq_num_dec_latch[2] ,
    \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/tx_hdr_seq_num_dec_latch[1] ,
    \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/tx_hdr_seq_num_dec_latch[0] ,
    \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/tx_lgood_empty ,
    \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/tx_lcrd_empty ,
    \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/send_hp_state[2] ,
    \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/send_hp_state[1] ,
    \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/send_hp_state[0] ,
    \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/send_lcmd_state[3] ,
    \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/send_lcmd_state[2] ,
    \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/send_lcmd_state[1] ,
    \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/send_lcmd_state[0] ,
    \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/tx_sel[2] ,
    \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/tx_sel[1] ,
    \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/tx_sel[0] ,
    \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/tx_lcrd_act ,
    \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/qc[7] ,
    \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/qc[6] ,
    \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/qc[5] ,
    \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/qc[4] ,
    \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/qc[3] ,
    \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/qc[2] ,
    \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/qc[1] ,
    \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/qc[0] ,
    \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/tx_lgood_act ,
    \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/res_state[2] ,
    \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/res_state[1] ,
    \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/res_state[0] ,
    \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/buf_out_dp_acked[2] ,
    \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/usb3_ep2_IN/buf_in_ready ,
    \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/usb3_ep2_IN/buf_in_commit ,
    \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/usb3_ep2_IN/buf_in_eob ,
    \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/usb3_ep2_IN/in_ep_rty ,
    \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/usb3_ep2_IN/buf_out_hasdata ,
    \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/usb3_ep2_IN/buf_out_eob ,
    \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/usb3_ep2_IN/buf_out_nump[4] ,
    \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/usb3_ep2_IN/buf_out_nump[3] ,
    \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/usb3_ep2_IN/buf_out_nump[2] ,
    \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/usb3_ep2_IN/buf_out_nump[1] ,
    \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/usb3_ep2_IN/buf_out_nump[0] ,
    \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/usb3_ep2_IN/buf_out_next_dp_ack_pt[3] ,
    \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/usb3_ep2_IN/buf_out_next_dp_ack_pt[2] ,
    \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/usb3_ep2_IN/buf_out_next_dp_ack_pt[1] ,
    \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/usb3_ep2_IN/buf_out_next_dp_ack_pt[0] ,
    \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/usb3_ep2_IN/buf_wt_ack_mem[15] ,
    \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/usb3_ep2_IN/buf_wt_ack_mem[14] ,
    \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/usb3_ep2_IN/buf_wt_ack_mem[13] ,
    \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/usb3_ep2_IN/buf_wt_ack_mem[12] ,
    \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/usb3_ep2_IN/buf_wt_ack_mem[11] ,
    \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/usb3_ep2_IN/buf_wt_ack_mem[10] ,
    \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/usb3_ep2_IN/buf_wt_ack_mem[9] ,
    \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/usb3_ep2_IN/buf_wt_ack_mem[8] ,
    \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/usb3_ep2_IN/buf_wt_ack_mem[7] ,
    \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/usb3_ep2_IN/buf_wt_ack_mem[6] ,
    \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/usb3_ep2_IN/buf_wt_ack_mem[5] ,
    \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/usb3_ep2_IN/buf_wt_ack_mem[4] ,
    \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/usb3_ep2_IN/buf_wt_ack_mem[3] ,
    \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/usb3_ep2_IN/buf_wt_ack_mem[2] ,
    \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/usb3_ep2_IN/buf_wt_ack_mem[1] ,
    \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/usb3_ep2_IN/buf_wt_ack_mem[0] ,
    \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/usb3_ep2_IN/buf_ready_mem[0] ,
    \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/usb3_ep2_IN/buf_ready_mem[1] ,
    \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/usb3_ep2_IN/buf_ready_mem[2] ,
    \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/usb3_ep2_IN/buf_ready_mem[3] ,
    \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/usb3_ep2_IN/buf_ready_mem[4] ,
    \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/usb3_ep2_IN/buf_ready_mem[5] ,
    \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/usb3_ep2_IN/buf_ready_mem[6] ,
    \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/usb3_ep2_IN/buf_ready_mem[7] ,
    \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/usb3_ep2_IN/buf_ready_mem[8] ,
    \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/usb3_ep2_IN/buf_ready_mem[9] ,
    \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/usb3_ep2_IN/buf_ready_mem[10] ,
    \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/usb3_ep2_IN/buf_ready_mem[11] ,
    \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/usb3_ep2_IN/buf_ready_mem[12] ,
    \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/usb3_ep2_IN/buf_ready_mem[13] ,
    \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/usb3_ep2_IN/buf_ready_mem[14] ,
    \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/usb3_ep2_IN/buf_ready_mem[15] ,
    \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/usb3_ep2_IN/buf_out_hasdata_mem[0] ,
    \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/usb3_ep2_IN/buf_out_hasdata_mem[1] ,
    \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/usb3_ep2_IN/buf_out_hasdata_mem[2] ,
    \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/usb3_ep2_IN/buf_out_hasdata_mem[3] ,
    \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/usb3_ep2_IN/buf_out_hasdata_mem[4] ,
    \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/usb3_ep2_IN/buf_out_hasdata_mem[5] ,
    \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/usb3_ep2_IN/buf_out_hasdata_mem[6] ,
    \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/usb3_ep2_IN/buf_out_hasdata_mem[7] ,
    \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/usb3_ep2_IN/buf_out_hasdata_mem[8] ,
    \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/usb3_ep2_IN/buf_out_hasdata_mem[9] ,
    \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/usb3_ep2_IN/buf_out_hasdata_mem[10] ,
    \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/usb3_ep2_IN/buf_out_hasdata_mem[11] ,
    \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/usb3_ep2_IN/buf_out_hasdata_mem[12] ,
    \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/usb3_ep2_IN/buf_out_hasdata_mem[13] ,
    \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/usb3_ep2_IN/buf_out_hasdata_mem[14] ,
    \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/usb3_ep2_IN/buf_out_hasdata_mem[15] ,
    \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/err_lbad_recv_latch ,
    \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/err_lbad_recv_latch_2 ,
    \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/usb3_ep2_IN/buf_out_pt[3] ,
    \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/usb3_ep2_IN/buf_out_pt[2] ,
    \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/usb3_ep2_IN/buf_out_pt[1] ,
    \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/usb3_ep2_IN/buf_out_pt[0] ,
    \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/usb3_ep2_IN/buf_in_pt[3] ,
    \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/usb3_ep2_IN/buf_in_pt[2] ,
    \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/usb3_ep2_IN/buf_in_pt[1] ,
    \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/usb3_ep2_IN/buf_in_pt[0] ,
    \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/usb3_ep2_IN/wt_ack_pt[3] ,
    \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/usb3_ep2_IN/wt_ack_pt[2] ,
    \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/usb3_ep2_IN/wt_ack_pt[1] ,
    \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/usb3_ep2_IN/wt_ack_pt[0] ,
    \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/tx_hp_act ,
    \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/err_hp_seq_latch ,
    \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/err_lgood_order_latch ,
    \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/tx_lgood_pop ,
    request_active,
    ep2_in_buf_data_commit,
    ep2_in_buf_eob,
    \UserLayer_top_inst/cam_active ,
    \dbg_ltssm_state[4] ,
    \dbg_ltssm_state[3] ,
    \dbg_ltssm_state[2] ,
    \dbg_ltssm_state[1] ,
    \dbg_ltssm_state[0] ,
    pclk,
    tms_pad_i,
    tck_pad_i,
    tdi_pad_i,
    tdo_pad_o
);

input \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/in_data[31] ;
input \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/in_data[30] ;
input \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/in_data[29] ;
input \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/in_data[28] ;
input \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/in_data[27] ;
input \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/in_data[26] ;
input \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/in_data[25] ;
input \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/in_data[24] ;
input \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/in_data[23] ;
input \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/in_data[22] ;
input \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/in_data[21] ;
input \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/in_data[20] ;
input \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/in_data[19] ;
input \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/in_data[18] ;
input \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/in_data[17] ;
input \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/in_data[16] ;
input \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/in_data[15] ;
input \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/in_data[14] ;
input \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/in_data[13] ;
input \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/in_data[12] ;
input \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/in_data[11] ;
input \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/in_data[10] ;
input \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/in_data[9] ;
input \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/in_data[8] ;
input \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/in_data[7] ;
input \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/in_data[6] ;
input \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/in_data[5] ;
input \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/in_data[4] ;
input \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/in_data[3] ;
input \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/in_data[2] ;
input \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/in_data[1] ;
input \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/in_data[0] ;
input \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/in_datak[3] ;
input \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/in_datak[2] ;
input \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/in_datak[1] ;
input \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/in_datak[0] ;
input \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/in_active ;
input \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/outp_data[31] ;
input \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/outp_data[30] ;
input \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/outp_data[29] ;
input \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/outp_data[28] ;
input \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/outp_data[27] ;
input \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/outp_data[26] ;
input \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/outp_data[25] ;
input \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/outp_data[24] ;
input \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/outp_data[23] ;
input \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/outp_data[22] ;
input \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/outp_data[21] ;
input \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/outp_data[20] ;
input \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/outp_data[19] ;
input \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/outp_data[18] ;
input \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/outp_data[17] ;
input \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/outp_data[16] ;
input \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/outp_data[15] ;
input \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/outp_data[14] ;
input \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/outp_data[13] ;
input \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/outp_data[12] ;
input \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/outp_data[11] ;
input \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/outp_data[10] ;
input \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/outp_data[9] ;
input \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/outp_data[8] ;
input \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/outp_data[7] ;
input \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/outp_data[6] ;
input \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/outp_data[5] ;
input \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/outp_data[4] ;
input \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/outp_data[3] ;
input \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/outp_data[2] ;
input \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/outp_data[1] ;
input \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/outp_data[0] ;
input \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/outp_datak[3] ;
input \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/outp_datak[2] ;
input \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/outp_datak[1] ;
input \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/outp_datak[0] ;
input \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/outp_active ;
input \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/out_stall ;
input \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/enter_u0_cnt[7] ;
input \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/enter_u0_cnt[6] ;
input \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/enter_u0_cnt[5] ;
input \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/enter_u0_cnt[4] ;
input \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/enter_u0_cnt[3] ;
input \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/enter_u0_cnt[2] ;
input \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/enter_u0_cnt[1] ;
input \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/enter_u0_cnt[0] ;
input \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/ltssm_exit_u0 ;
input \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/ltssm_current_state[4] ;
input \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/ltssm_current_state[3] ;
input \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/ltssm_current_state[2] ;
input \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/ltssm_current_state[1] ;
input \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/ltssm_current_state[0] ;
input \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/queue_send_u0_adv ;
input \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/queue_send_u0_portcap ;
input \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/link_cmd_det ;
input \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/send_port_cfg_resp ;
input \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/remote_rx_cred_count[2] ;
input \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/remote_rx_cred_count[1] ;
input \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/remote_rx_cred_count[0] ;
input \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/tx_cred_idx[1] ;
input \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/tx_cred_idx[0] ;
input \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/send_port_cfg_resp_ack ;
input \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/ack_tx_hdr_seq_num[2] ;
input \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/ack_tx_hdr_seq_num[1] ;
input \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/ack_tx_hdr_seq_num[0] ;
input \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/rx_hdr_seq_num[2] ;
input \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/rx_hdr_seq_num[1] ;
input \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/rx_hdr_seq_num[0] ;
input \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/ltssm_enter_u0_by_polling ;
input \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/in_link_command_act ;
input \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/in_link_command_crc_good ;
input \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/in_link_command_latch_act ;
input \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/recv_u0_adv ;
input \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/err_lgood_order ;
input \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/err_lcrd_mismatch ;
input \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/err_lbad_recv ;
input \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/hp_det ;
input \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/in_header_act ;
input \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/hp_crc_good ;
input \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/err_hp_seq ;
input \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/err_lbad ;
input \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/local_rx_cred_count[2] ;
input \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/local_rx_cred_count[1] ;
input \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/local_rx_cred_count[0] ;
input \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/rx_dph ;
input \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/rx_dph_eob ;
input \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/rx_dph_setup ;
input \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/rx_dph_pktpend ;
input \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/rx_dph_endp[3] ;
input \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/rx_dph_endp[2] ;
input \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/rx_dph_endp[1] ;
input \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/rx_dph_endp[0] ;
input \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/rx_dph_seq[4] ;
input \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/rx_dph_seq[3] ;
input \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/rx_dph_seq[2] ;
input \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/rx_dph_seq[1] ;
input \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/rx_dph_seq[0] ;
input \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/rx_dph_len[15] ;
input \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/rx_dph_len[14] ;
input \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/rx_dph_len[13] ;
input \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/rx_dph_len[12] ;
input \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/rx_dph_len[11] ;
input \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/rx_dph_len[10] ;
input \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/rx_dph_len[9] ;
input \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/rx_dph_len[8] ;
input \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/rx_dph_len[7] ;
input \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/rx_dph_len[6] ;
input \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/rx_dph_len[5] ;
input \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/rx_dph_len[4] ;
input \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/rx_dph_len[3] ;
input \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/rx_dph_len[2] ;
input \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/rx_dph_len[1] ;
input \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/rx_dph_len[0] ;
input \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/rx_tp_subtype[3] ;
input \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/rx_tp_subtype[2] ;
input \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/rx_tp_subtype[1] ;
input \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/rx_tp_subtype[0] ;
input \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/rx_tp_endp[3] ;
input \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/rx_tp_endp[2] ;
input \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/rx_tp_endp[1] ;
input \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/rx_tp_endp[0] ;
input \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/rx_tp_nump[4] ;
input \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/rx_tp_nump[3] ;
input \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/rx_tp_nump[2] ;
input \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/rx_tp_nump[1] ;
input \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/rx_tp_nump[0] ;
input \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/rx_tp_seq[4] ;
input \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/rx_tp_seq[3] ;
input \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/rx_tp_seq[2] ;
input \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/rx_tp_seq[1] ;
input \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/rx_tp_seq[0] ;
input \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/rx_tp_stream[15] ;
input \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/rx_tp_stream[14] ;
input \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/rx_tp_stream[13] ;
input \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/rx_tp_stream[12] ;
input \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/rx_tp_stream[11] ;
input \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/rx_tp_stream[10] ;
input \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/rx_tp_stream[9] ;
input \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/rx_tp_stream[8] ;
input \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/rx_tp_stream[7] ;
input \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/rx_tp_stream[6] ;
input \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/rx_tp_stream[5] ;
input \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/rx_tp_stream[4] ;
input \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/rx_tp_stream[3] ;
input \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/rx_tp_stream[2] ;
input \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/rx_tp_stream[1] ;
input \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/rx_tp_stream[0] ;
input \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/rx_tp ;
input \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/rx_tp_retry ;
input \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/rx_tp_pktpend ;
input \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/tx_tp_a_subtype[3] ;
input \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/tx_tp_a_subtype[2] ;
input \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/tx_tp_a_subtype[1] ;
input \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/tx_tp_a_subtype[0] ;
input \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/tx_tp_a_endp[3] ;
input \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/tx_tp_a_endp[2] ;
input \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/tx_tp_a_endp[1] ;
input \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/tx_tp_a_endp[0] ;
input \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/tx_tp_a ;
input \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/tx_tp_a_dir ;
input \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/tx_tp_a_nump[4] ;
input \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/tx_tp_a_nump[3] ;
input \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/tx_tp_a_nump[2] ;
input \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/tx_tp_a_nump[1] ;
input \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/tx_tp_a_nump[0] ;
input \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/tx_tp_a_seq[4] ;
input \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/tx_tp_a_seq[3] ;
input \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/tx_tp_a_seq[2] ;
input \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/tx_tp_a_seq[1] ;
input \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/tx_tp_a_seq[0] ;
input \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/tx_tp_a_stream[15] ;
input \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/tx_tp_a_stream[14] ;
input \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/tx_tp_a_stream[13] ;
input \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/tx_tp_a_stream[12] ;
input \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/tx_tp_a_stream[11] ;
input \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/tx_tp_a_stream[10] ;
input \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/tx_tp_a_stream[9] ;
input \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/tx_tp_a_stream[8] ;
input \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/tx_tp_a_stream[7] ;
input \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/tx_tp_a_stream[6] ;
input \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/tx_tp_a_stream[5] ;
input \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/tx_tp_a_stream[4] ;
input \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/tx_tp_a_stream[3] ;
input \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/tx_tp_a_stream[2] ;
input \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/tx_tp_a_stream[1] ;
input \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/tx_tp_a_stream[0] ;
input \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/tx_tp_a_retry ;
input \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/tx_tp_b_subtype[3] ;
input \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/tx_tp_b_subtype[2] ;
input \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/tx_tp_b_subtype[1] ;
input \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/tx_tp_b_subtype[0] ;
input \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/tx_tp_b_endp[3] ;
input \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/tx_tp_b_endp[2] ;
input \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/tx_tp_b_endp[1] ;
input \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/tx_tp_b_endp[0] ;
input \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/tx_tp_b ;
input \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/tx_tp_b_retry ;
input \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/tx_tp_b_nump[4] ;
input \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/tx_tp_b_nump[3] ;
input \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/tx_tp_b_nump[2] ;
input \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/tx_tp_b_nump[1] ;
input \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/tx_tp_b_nump[0] ;
input \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/tx_tp_c_subtype[3] ;
input \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/tx_tp_c_subtype[2] ;
input \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/tx_tp_c_subtype[1] ;
input \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/tx_tp_c_subtype[0] ;
input \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/tx_tp_c_endp[3] ;
input \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/tx_tp_c_endp[2] ;
input \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/tx_tp_c_endp[1] ;
input \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/tx_tp_c_endp[0] ;
input \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/tx_tp_c ;
input \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/tx_tp_c_retry ;
input \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/tx_tp_c_nump[4] ;
input \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/tx_tp_c_nump[3] ;
input \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/tx_tp_c_nump[2] ;
input \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/tx_tp_c_nump[1] ;
input \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/tx_tp_c_nump[0] ;
input \UserLayer_top_inst/DataTransfer_inst/ep1_in_buf_ready ;
input \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/iu3ep0/req_cnt[7] ;
input \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/iu3ep0/req_cnt[6] ;
input \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/iu3ep0/req_cnt[5] ;
input \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/iu3ep0/req_cnt[4] ;
input \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/iu3ep0/req_cnt[3] ;
input \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/iu3ep0/req_cnt[2] ;
input \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/iu3ep0/req_cnt[1] ;
input \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/iu3ep0/req_cnt[0] ;
input \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/host_requests_data ;
input \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/host_requests_endpt[3] ;
input \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/host_requests_endpt[2] ;
input \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/host_requests_endpt[1] ;
input \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/host_requests_endpt[0] ;
input \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/rx_dpp_start ;
input \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/rx_dpp_done ;
input \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/rx_dpp_crcgood ;
input \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/err_missed_dpp_start ;
input \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/err_missed_dpp_done ;
input \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/tx_dph ;
input \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/tx_dph_eob ;
input \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/tx_dph_dir ;
input \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/tx_dph_endp[3] ;
input \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/tx_dph_endp[2] ;
input \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/tx_dph_endp[1] ;
input \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/tx_dph_endp[0] ;
input \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/tx_dph_seq[4] ;
input \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/tx_dph_seq[3] ;
input \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/tx_dph_seq[2] ;
input \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/tx_dph_seq[1] ;
input \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/tx_dph_seq[0] ;
input \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/tx_dph_len[15] ;
input \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/tx_dph_len[14] ;
input \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/tx_dph_len[13] ;
input \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/tx_dph_len[12] ;
input \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/tx_dph_len[11] ;
input \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/tx_dph_len[10] ;
input \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/tx_dph_len[9] ;
input \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/tx_dph_len[8] ;
input \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/tx_dph_len[7] ;
input \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/tx_dph_len[6] ;
input \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/tx_dph_len[5] ;
input \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/tx_dph_len[4] ;
input \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/tx_dph_len[3] ;
input \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/tx_dph_len[2] ;
input \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/tx_dph_len[1] ;
input \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/tx_dph_len[0] ;
input \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/tx_dpp_ack ;
input \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/tx_dpp_done ;
input \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/ep2_buf_out_nump[4] ;
input \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/ep2_buf_out_nump[3] ;
input \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/ep2_buf_out_nump[2] ;
input \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/ep2_buf_out_nump[1] ;
input \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/ep2_buf_out_nump[0] ;
input \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/burst_in_act ;
input \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/burst_in_stop ;
input \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/do_send_dpp ;
input \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/do_send_dpp_ack ;
input \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/do_send_dpp_eob ;
input \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/crc_hprx_out[15] ;
input \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/crc_hprx_out[14] ;
input \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/crc_hprx_out[13] ;
input \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/crc_hprx_out[12] ;
input \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/crc_hprx_out[11] ;
input \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/crc_hprx_out[10] ;
input \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/crc_hprx_out[9] ;
input \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/crc_hprx_out[8] ;
input \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/crc_hprx_out[7] ;
input \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/crc_hprx_out[6] ;
input \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/crc_hprx_out[5] ;
input \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/crc_hprx_out[4] ;
input \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/crc_hprx_out[3] ;
input \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/crc_hprx_out[2] ;
input \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/crc_hprx_out[1] ;
input \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/crc_hprx_out[0] ;
input \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/crc_hprx_rst ;
input \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/crc_hprx_en ;
input \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/crc_hprx_in[31] ;
input \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/crc_hprx_in[30] ;
input \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/crc_hprx_in[29] ;
input \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/crc_hprx_in[28] ;
input \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/crc_hprx_in[27] ;
input \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/crc_hprx_in[26] ;
input \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/crc_hprx_in[25] ;
input \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/crc_hprx_in[24] ;
input \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/crc_hprx_in[23] ;
input \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/crc_hprx_in[22] ;
input \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/crc_hprx_in[21] ;
input \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/crc_hprx_in[20] ;
input \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/crc_hprx_in[19] ;
input \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/crc_hprx_in[18] ;
input \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/crc_hprx_in[17] ;
input \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/crc_hprx_in[16] ;
input \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/crc_hprx_in[15] ;
input \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/crc_hprx_in[14] ;
input \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/crc_hprx_in[13] ;
input \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/crc_hprx_in[12] ;
input \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/crc_hprx_in[11] ;
input \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/crc_hprx_in[10] ;
input \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/crc_hprx_in[9] ;
input \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/crc_hprx_in[8] ;
input \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/crc_hprx_in[7] ;
input \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/crc_hprx_in[6] ;
input \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/crc_hprx_in[5] ;
input \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/crc_hprx_in[4] ;
input \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/crc_hprx_in[3] ;
input \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/crc_hprx_in[2] ;
input \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/crc_hprx_in[1] ;
input \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/crc_hprx_in[0] ;
input \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/crc_cw3_out[4] ;
input \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/crc_cw3_out[3] ;
input \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/crc_cw3_out[2] ;
input \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/crc_cw3_out[1] ;
input \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/crc_cw3_out[0] ;
input \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/in_header_cw[15] ;
input \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/in_header_cw[14] ;
input \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/in_header_cw[13] ;
input \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/in_header_cw[12] ;
input \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/in_header_cw[11] ;
input \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/in_header_cw[10] ;
input \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/in_header_cw[9] ;
input \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/in_header_cw[8] ;
input \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/in_header_cw[7] ;
input \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/in_header_cw[6] ;
input \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/in_header_cw[5] ;
input \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/in_header_cw[4] ;
input \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/in_header_cw[3] ;
input \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/in_header_cw[2] ;
input \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/in_header_cw[1] ;
input \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/in_header_cw[0] ;
input \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/in_link_command[10] ;
input \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/in_link_command[9] ;
input \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/in_link_command[8] ;
input \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/in_link_command[7] ;
input \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/in_link_command[6] ;
input \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/in_link_command[5] ;
input \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/in_link_command[4] ;
input \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/in_link_command[3] ;
input \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/in_link_command[2] ;
input \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/in_link_command[1] ;
input \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/in_link_command[0] ;
input \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/crc_cw1_out[4] ;
input \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/crc_cw1_out[3] ;
input \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/crc_cw1_out[2] ;
input \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/crc_cw1_out[1] ;
input \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/crc_cw1_out[0] ;
input \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/in_link_command[31] ;
input \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/in_link_command[30] ;
input \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/in_link_command[29] ;
input \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/in_link_command[28] ;
input \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/in_link_command[27] ;
input \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/in_link_command[26] ;
input \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/in_link_command[25] ;
input \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/in_link_command[24] ;
input \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/in_link_command[23] ;
input \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/in_link_command[22] ;
input \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/in_link_command[21] ;
input \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/in_link_command[20] ;
input \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/in_link_command[19] ;
input \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/in_link_command[18] ;
input \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/in_link_command[17] ;
input \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/in_link_command[16] ;
input \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/crc_cw2_out[4] ;
input \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/crc_cw2_out[3] ;
input \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/crc_cw2_out[2] ;
input \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/crc_cw2_out[1] ;
input \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/crc_cw2_out[0] ;
input \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/in_link_command[15] ;
input \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/in_link_command[14] ;
input \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/in_link_command[13] ;
input \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/in_link_command[12] ;
input \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/in_link_command[11] ;
input \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/err_lbad_reg ;
input \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/rx_hdr_seq_num_reg[2] ;
input \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/rx_hdr_seq_num_reg[1] ;
input \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/rx_hdr_seq_num_reg[0] ;
input \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/link_err ;
input \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/tx_lbad_pop ;
input \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/tx_lbad_q[10] ;
input \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/tx_lbad_q[9] ;
input \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/tx_lbad_q[8] ;
input \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/tx_lbad_q[7] ;
input \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/tx_lbad_q[6] ;
input \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/tx_lbad_q[5] ;
input \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/tx_lbad_q[4] ;
input \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/tx_lbad_q[3] ;
input \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/tx_lbad_q[2] ;
input \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/tx_lbad_q[1] ;
input \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/tx_lbad_q[0] ;
input \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/tx_lbad_empty ;
input \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/tx_lbad_act ;
input \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/wait_retry ;
input \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/rx_retry ;
input \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/hp_valid_k_cnt[2] ;
input \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/hp_valid_k_cnt[1] ;
input \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/hp_valid_k_cnt[0] ;
input \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/hp_valid_k[3] ;
input \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/hp_valid_k[2] ;
input \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/hp_valid_k[1] ;
input \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/hp_valid_k[0] ;
input \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/queue_state[2] ;
input \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/queue_state[1] ;
input \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/queue_state[0] ;
input \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/send_dpp_state[3] ;
input \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/send_dpp_state[2] ;
input \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/send_dpp_state[1] ;
input \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/send_dpp_state[0] ;
input \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/tx_link_busy ;
input \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/tx_lcmd_req ;
input \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/tx_hp_req ;
input \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/ltssm_state[4] ;
input \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/ltssm_state[3] ;
input \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/ltssm_state[2] ;
input \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/ltssm_state[1] ;
input \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/ltssm_state[0] ;
input \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/reset_n ;
input \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/ltssm_go_recovery ;
input \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/res_mem_wr_en ;
input \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/res_mem_wr_dat[35] ;
input \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/res_mem_wr_dat[34] ;
input \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/res_mem_wr_dat[33] ;
input \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/res_mem_wr_dat[32] ;
input \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/res_mem_wr_dat[31] ;
input \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/res_mem_wr_dat[30] ;
input \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/res_mem_wr_dat[29] ;
input \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/res_mem_wr_dat[28] ;
input \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/res_mem_wr_dat[27] ;
input \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/res_mem_wr_dat[26] ;
input \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/res_mem_wr_dat[25] ;
input \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/res_mem_wr_dat[24] ;
input \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/res_mem_wr_dat[23] ;
input \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/res_mem_wr_dat[22] ;
input \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/res_mem_wr_dat[21] ;
input \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/res_mem_wr_dat[20] ;
input \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/res_mem_wr_dat[19] ;
input \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/res_mem_wr_dat[18] ;
input \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/res_mem_wr_dat[17] ;
input \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/res_mem_wr_dat[16] ;
input \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/res_mem_wr_dat[15] ;
input \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/res_mem_wr_dat[14] ;
input \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/res_mem_wr_dat[13] ;
input \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/res_mem_wr_dat[12] ;
input \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/res_mem_wr_dat[11] ;
input \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/res_mem_wr_dat[10] ;
input \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/res_mem_wr_dat[9] ;
input \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/res_mem_wr_dat[8] ;
input \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/res_mem_wr_dat[7] ;
input \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/res_mem_wr_dat[6] ;
input \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/res_mem_wr_dat[5] ;
input \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/res_mem_wr_dat[4] ;
input \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/res_mem_wr_dat[3] ;
input \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/res_mem_wr_dat[2] ;
input \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/res_mem_wr_dat[1] ;
input \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/res_mem_wr_dat[0] ;
input \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/res_mem_wr_addr[10] ;
input \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/res_mem_wr_addr[9] ;
input \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/res_mem_wr_addr[8] ;
input \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/res_mem_wr_addr[7] ;
input \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/res_mem_wr_addr[6] ;
input \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/res_mem_wr_addr[5] ;
input \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/res_mem_wr_addr[4] ;
input \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/res_mem_wr_addr[3] ;
input \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/res_mem_wr_addr[2] ;
input \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/res_mem_wr_addr[1] ;
input \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/res_mem_wr_addr[0] ;
input \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/res_mem_wr_pt[1] ;
input \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/res_mem_wr_pt[0] ;
input \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/resend_hp_act ;
input \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/tx_hdr_seq_num_dec[2] ;
input \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/tx_hdr_seq_num_dec[1] ;
input \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/tx_hdr_seq_num_dec[0] ;
input \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/resend_hp_num[4] ;
input \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/resend_hp_num[3] ;
input \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/resend_hp_num[2] ;
input \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/resend_hp_num[1] ;
input \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/resend_hp_num[0] ;
input \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/res_mem_rd_pt[1] ;
input \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/res_mem_rd_pt[0] ;
input \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/res_mem_rd_addr[10] ;
input \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/res_mem_rd_addr[9] ;
input \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/res_mem_rd_addr[8] ;
input \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/res_mem_rd_addr[7] ;
input \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/res_mem_rd_addr[6] ;
input \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/res_mem_rd_addr[5] ;
input \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/res_mem_rd_addr[4] ;
input \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/res_mem_rd_addr[3] ;
input \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/res_mem_rd_addr[2] ;
input \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/res_mem_rd_addr[1] ;
input \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/res_mem_rd_addr[0] ;
input \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/res_mem_rd_en ;
input \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/tx_res_req ;
input \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/tx_res_req_ack ;
input \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/res_mem_rd_dat[35] ;
input \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/res_mem_rd_dat[34] ;
input \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/res_mem_rd_dat[33] ;
input \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/res_mem_rd_dat[32] ;
input \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/res_mem_rd_dat[31] ;
input \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/res_mem_rd_dat[30] ;
input \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/res_mem_rd_dat[29] ;
input \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/res_mem_rd_dat[28] ;
input \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/res_mem_rd_dat[27] ;
input \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/res_mem_rd_dat[26] ;
input \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/res_mem_rd_dat[25] ;
input \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/res_mem_rd_dat[24] ;
input \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/res_mem_rd_dat[23] ;
input \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/res_mem_rd_dat[22] ;
input \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/res_mem_rd_dat[21] ;
input \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/res_mem_rd_dat[20] ;
input \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/res_mem_rd_dat[19] ;
input \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/res_mem_rd_dat[18] ;
input \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/res_mem_rd_dat[17] ;
input \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/res_mem_rd_dat[16] ;
input \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/res_mem_rd_dat[15] ;
input \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/res_mem_rd_dat[14] ;
input \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/res_mem_rd_dat[13] ;
input \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/res_mem_rd_dat[12] ;
input \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/res_mem_rd_dat[11] ;
input \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/res_mem_rd_dat[10] ;
input \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/res_mem_rd_dat[9] ;
input \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/res_mem_rd_dat[8] ;
input \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/res_mem_rd_dat[7] ;
input \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/res_mem_rd_dat[6] ;
input \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/res_mem_rd_dat[5] ;
input \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/res_mem_rd_dat[4] ;
input \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/res_mem_rd_dat[3] ;
input \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/res_mem_rd_dat[2] ;
input \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/res_mem_rd_dat[1] ;
input \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/res_mem_rd_dat[0] ;
input \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/res_mem_rd_dat_val ;
input \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/out_data_5[31] ;
input \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/out_data_5[30] ;
input \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/out_data_5[29] ;
input \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/out_data_5[28] ;
input \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/out_data_5[27] ;
input \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/out_data_5[26] ;
input \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/out_data_5[25] ;
input \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/out_data_5[24] ;
input \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/out_data_5[23] ;
input \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/out_data_5[22] ;
input \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/out_data_5[21] ;
input \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/out_data_5[20] ;
input \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/out_data_5[19] ;
input \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/out_data_5[18] ;
input \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/out_data_5[17] ;
input \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/out_data_5[16] ;
input \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/out_data_5[15] ;
input \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/out_data_5[14] ;
input \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/out_data_5[13] ;
input \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/out_data_5[12] ;
input \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/out_data_5[11] ;
input \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/out_data_5[10] ;
input \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/out_data_5[9] ;
input \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/out_data_5[8] ;
input \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/out_data_5[7] ;
input \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/out_data_5[6] ;
input \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/out_data_5[5] ;
input \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/out_data_5[4] ;
input \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/out_data_5[3] ;
input \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/out_data_5[2] ;
input \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/out_data_5[1] ;
input \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/out_data_5[0] ;
input \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/out_datak_5[3] ;
input \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/out_datak_5[2] ;
input \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/out_datak_5[1] ;
input \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/out_datak_5[0] ;
input \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/out_active_5 ;
input \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/tx_hdr_seq_num_dec_latch[2] ;
input \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/tx_hdr_seq_num_dec_latch[1] ;
input \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/tx_hdr_seq_num_dec_latch[0] ;
input \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/tx_lgood_empty ;
input \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/tx_lcrd_empty ;
input \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/send_hp_state[2] ;
input \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/send_hp_state[1] ;
input \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/send_hp_state[0] ;
input \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/send_lcmd_state[3] ;
input \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/send_lcmd_state[2] ;
input \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/send_lcmd_state[1] ;
input \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/send_lcmd_state[0] ;
input \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/tx_sel[2] ;
input \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/tx_sel[1] ;
input \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/tx_sel[0] ;
input \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/tx_lcrd_act ;
input \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/qc[7] ;
input \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/qc[6] ;
input \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/qc[5] ;
input \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/qc[4] ;
input \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/qc[3] ;
input \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/qc[2] ;
input \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/qc[1] ;
input \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/qc[0] ;
input \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/tx_lgood_act ;
input \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/res_state[2] ;
input \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/res_state[1] ;
input \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/res_state[0] ;
input \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/buf_out_dp_acked[2] ;
input \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/usb3_ep2_IN/buf_in_ready ;
input \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/usb3_ep2_IN/buf_in_commit ;
input \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/usb3_ep2_IN/buf_in_eob ;
input \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/usb3_ep2_IN/in_ep_rty ;
input \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/usb3_ep2_IN/buf_out_hasdata ;
input \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/usb3_ep2_IN/buf_out_eob ;
input \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/usb3_ep2_IN/buf_out_nump[4] ;
input \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/usb3_ep2_IN/buf_out_nump[3] ;
input \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/usb3_ep2_IN/buf_out_nump[2] ;
input \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/usb3_ep2_IN/buf_out_nump[1] ;
input \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/usb3_ep2_IN/buf_out_nump[0] ;
input \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/usb3_ep2_IN/buf_out_next_dp_ack_pt[3] ;
input \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/usb3_ep2_IN/buf_out_next_dp_ack_pt[2] ;
input \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/usb3_ep2_IN/buf_out_next_dp_ack_pt[1] ;
input \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/usb3_ep2_IN/buf_out_next_dp_ack_pt[0] ;
input \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/usb3_ep2_IN/buf_wt_ack_mem[15] ;
input \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/usb3_ep2_IN/buf_wt_ack_mem[14] ;
input \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/usb3_ep2_IN/buf_wt_ack_mem[13] ;
input \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/usb3_ep2_IN/buf_wt_ack_mem[12] ;
input \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/usb3_ep2_IN/buf_wt_ack_mem[11] ;
input \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/usb3_ep2_IN/buf_wt_ack_mem[10] ;
input \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/usb3_ep2_IN/buf_wt_ack_mem[9] ;
input \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/usb3_ep2_IN/buf_wt_ack_mem[8] ;
input \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/usb3_ep2_IN/buf_wt_ack_mem[7] ;
input \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/usb3_ep2_IN/buf_wt_ack_mem[6] ;
input \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/usb3_ep2_IN/buf_wt_ack_mem[5] ;
input \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/usb3_ep2_IN/buf_wt_ack_mem[4] ;
input \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/usb3_ep2_IN/buf_wt_ack_mem[3] ;
input \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/usb3_ep2_IN/buf_wt_ack_mem[2] ;
input \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/usb3_ep2_IN/buf_wt_ack_mem[1] ;
input \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/usb3_ep2_IN/buf_wt_ack_mem[0] ;
input \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/usb3_ep2_IN/buf_ready_mem[0] ;
input \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/usb3_ep2_IN/buf_ready_mem[1] ;
input \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/usb3_ep2_IN/buf_ready_mem[2] ;
input \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/usb3_ep2_IN/buf_ready_mem[3] ;
input \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/usb3_ep2_IN/buf_ready_mem[4] ;
input \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/usb3_ep2_IN/buf_ready_mem[5] ;
input \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/usb3_ep2_IN/buf_ready_mem[6] ;
input \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/usb3_ep2_IN/buf_ready_mem[7] ;
input \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/usb3_ep2_IN/buf_ready_mem[8] ;
input \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/usb3_ep2_IN/buf_ready_mem[9] ;
input \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/usb3_ep2_IN/buf_ready_mem[10] ;
input \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/usb3_ep2_IN/buf_ready_mem[11] ;
input \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/usb3_ep2_IN/buf_ready_mem[12] ;
input \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/usb3_ep2_IN/buf_ready_mem[13] ;
input \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/usb3_ep2_IN/buf_ready_mem[14] ;
input \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/usb3_ep2_IN/buf_ready_mem[15] ;
input \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/usb3_ep2_IN/buf_out_hasdata_mem[0] ;
input \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/usb3_ep2_IN/buf_out_hasdata_mem[1] ;
input \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/usb3_ep2_IN/buf_out_hasdata_mem[2] ;
input \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/usb3_ep2_IN/buf_out_hasdata_mem[3] ;
input \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/usb3_ep2_IN/buf_out_hasdata_mem[4] ;
input \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/usb3_ep2_IN/buf_out_hasdata_mem[5] ;
input \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/usb3_ep2_IN/buf_out_hasdata_mem[6] ;
input \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/usb3_ep2_IN/buf_out_hasdata_mem[7] ;
input \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/usb3_ep2_IN/buf_out_hasdata_mem[8] ;
input \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/usb3_ep2_IN/buf_out_hasdata_mem[9] ;
input \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/usb3_ep2_IN/buf_out_hasdata_mem[10] ;
input \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/usb3_ep2_IN/buf_out_hasdata_mem[11] ;
input \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/usb3_ep2_IN/buf_out_hasdata_mem[12] ;
input \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/usb3_ep2_IN/buf_out_hasdata_mem[13] ;
input \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/usb3_ep2_IN/buf_out_hasdata_mem[14] ;
input \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/usb3_ep2_IN/buf_out_hasdata_mem[15] ;
input \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/err_lbad_recv_latch ;
input \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/err_lbad_recv_latch_2 ;
input \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/usb3_ep2_IN/buf_out_pt[3] ;
input \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/usb3_ep2_IN/buf_out_pt[2] ;
input \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/usb3_ep2_IN/buf_out_pt[1] ;
input \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/usb3_ep2_IN/buf_out_pt[0] ;
input \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/usb3_ep2_IN/buf_in_pt[3] ;
input \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/usb3_ep2_IN/buf_in_pt[2] ;
input \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/usb3_ep2_IN/buf_in_pt[1] ;
input \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/usb3_ep2_IN/buf_in_pt[0] ;
input \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/usb3_ep2_IN/wt_ack_pt[3] ;
input \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/usb3_ep2_IN/wt_ack_pt[2] ;
input \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/usb3_ep2_IN/wt_ack_pt[1] ;
input \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/usb3_ep2_IN/wt_ack_pt[0] ;
input \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/tx_hp_act ;
input \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/err_hp_seq_latch ;
input \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/err_lgood_order_latch ;
input \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/tx_lgood_pop ;
input request_active;
input ep2_in_buf_data_commit;
input ep2_in_buf_eob;
input \UserLayer_top_inst/cam_active ;
input \dbg_ltssm_state[4] ;
input \dbg_ltssm_state[3] ;
input \dbg_ltssm_state[2] ;
input \dbg_ltssm_state[1] ;
input \dbg_ltssm_state[0] ;
input pclk;
input tms_pad_i;
input tck_pad_i;
input tdi_pad_i;
output tdo_pad_o;

wire \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/in_data[31] ;
wire \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/in_data[30] ;
wire \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/in_data[29] ;
wire \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/in_data[28] ;
wire \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/in_data[27] ;
wire \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/in_data[26] ;
wire \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/in_data[25] ;
wire \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/in_data[24] ;
wire \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/in_data[23] ;
wire \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/in_data[22] ;
wire \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/in_data[21] ;
wire \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/in_data[20] ;
wire \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/in_data[19] ;
wire \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/in_data[18] ;
wire \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/in_data[17] ;
wire \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/in_data[16] ;
wire \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/in_data[15] ;
wire \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/in_data[14] ;
wire \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/in_data[13] ;
wire \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/in_data[12] ;
wire \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/in_data[11] ;
wire \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/in_data[10] ;
wire \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/in_data[9] ;
wire \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/in_data[8] ;
wire \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/in_data[7] ;
wire \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/in_data[6] ;
wire \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/in_data[5] ;
wire \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/in_data[4] ;
wire \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/in_data[3] ;
wire \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/in_data[2] ;
wire \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/in_data[1] ;
wire \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/in_data[0] ;
wire \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/in_datak[3] ;
wire \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/in_datak[2] ;
wire \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/in_datak[1] ;
wire \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/in_datak[0] ;
wire \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/in_active ;
wire \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/outp_data[31] ;
wire \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/outp_data[30] ;
wire \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/outp_data[29] ;
wire \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/outp_data[28] ;
wire \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/outp_data[27] ;
wire \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/outp_data[26] ;
wire \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/outp_data[25] ;
wire \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/outp_data[24] ;
wire \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/outp_data[23] ;
wire \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/outp_data[22] ;
wire \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/outp_data[21] ;
wire \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/outp_data[20] ;
wire \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/outp_data[19] ;
wire \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/outp_data[18] ;
wire \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/outp_data[17] ;
wire \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/outp_data[16] ;
wire \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/outp_data[15] ;
wire \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/outp_data[14] ;
wire \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/outp_data[13] ;
wire \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/outp_data[12] ;
wire \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/outp_data[11] ;
wire \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/outp_data[10] ;
wire \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/outp_data[9] ;
wire \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/outp_data[8] ;
wire \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/outp_data[7] ;
wire \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/outp_data[6] ;
wire \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/outp_data[5] ;
wire \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/outp_data[4] ;
wire \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/outp_data[3] ;
wire \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/outp_data[2] ;
wire \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/outp_data[1] ;
wire \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/outp_data[0] ;
wire \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/outp_datak[3] ;
wire \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/outp_datak[2] ;
wire \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/outp_datak[1] ;
wire \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/outp_datak[0] ;
wire \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/outp_active ;
wire \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/out_stall ;
wire \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/enter_u0_cnt[7] ;
wire \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/enter_u0_cnt[6] ;
wire \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/enter_u0_cnt[5] ;
wire \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/enter_u0_cnt[4] ;
wire \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/enter_u0_cnt[3] ;
wire \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/enter_u0_cnt[2] ;
wire \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/enter_u0_cnt[1] ;
wire \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/enter_u0_cnt[0] ;
wire \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/ltssm_exit_u0 ;
wire \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/ltssm_current_state[4] ;
wire \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/ltssm_current_state[3] ;
wire \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/ltssm_current_state[2] ;
wire \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/ltssm_current_state[1] ;
wire \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/ltssm_current_state[0] ;
wire \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/queue_send_u0_adv ;
wire \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/queue_send_u0_portcap ;
wire \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/link_cmd_det ;
wire \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/send_port_cfg_resp ;
wire \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/remote_rx_cred_count[2] ;
wire \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/remote_rx_cred_count[1] ;
wire \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/remote_rx_cred_count[0] ;
wire \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/tx_cred_idx[1] ;
wire \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/tx_cred_idx[0] ;
wire \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/send_port_cfg_resp_ack ;
wire \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/ack_tx_hdr_seq_num[2] ;
wire \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/ack_tx_hdr_seq_num[1] ;
wire \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/ack_tx_hdr_seq_num[0] ;
wire \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/rx_hdr_seq_num[2] ;
wire \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/rx_hdr_seq_num[1] ;
wire \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/rx_hdr_seq_num[0] ;
wire \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/ltssm_enter_u0_by_polling ;
wire \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/in_link_command_act ;
wire \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/in_link_command_crc_good ;
wire \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/in_link_command_latch_act ;
wire \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/recv_u0_adv ;
wire \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/err_lgood_order ;
wire \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/err_lcrd_mismatch ;
wire \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/err_lbad_recv ;
wire \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/hp_det ;
wire \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/in_header_act ;
wire \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/hp_crc_good ;
wire \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/err_hp_seq ;
wire \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/err_lbad ;
wire \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/local_rx_cred_count[2] ;
wire \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/local_rx_cred_count[1] ;
wire \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/local_rx_cred_count[0] ;
wire \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/rx_dph ;
wire \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/rx_dph_eob ;
wire \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/rx_dph_setup ;
wire \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/rx_dph_pktpend ;
wire \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/rx_dph_endp[3] ;
wire \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/rx_dph_endp[2] ;
wire \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/rx_dph_endp[1] ;
wire \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/rx_dph_endp[0] ;
wire \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/rx_dph_seq[4] ;
wire \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/rx_dph_seq[3] ;
wire \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/rx_dph_seq[2] ;
wire \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/rx_dph_seq[1] ;
wire \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/rx_dph_seq[0] ;
wire \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/rx_dph_len[15] ;
wire \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/rx_dph_len[14] ;
wire \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/rx_dph_len[13] ;
wire \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/rx_dph_len[12] ;
wire \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/rx_dph_len[11] ;
wire \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/rx_dph_len[10] ;
wire \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/rx_dph_len[9] ;
wire \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/rx_dph_len[8] ;
wire \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/rx_dph_len[7] ;
wire \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/rx_dph_len[6] ;
wire \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/rx_dph_len[5] ;
wire \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/rx_dph_len[4] ;
wire \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/rx_dph_len[3] ;
wire \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/rx_dph_len[2] ;
wire \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/rx_dph_len[1] ;
wire \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/rx_dph_len[0] ;
wire \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/rx_tp_subtype[3] ;
wire \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/rx_tp_subtype[2] ;
wire \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/rx_tp_subtype[1] ;
wire \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/rx_tp_subtype[0] ;
wire \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/rx_tp_endp[3] ;
wire \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/rx_tp_endp[2] ;
wire \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/rx_tp_endp[1] ;
wire \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/rx_tp_endp[0] ;
wire \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/rx_tp_nump[4] ;
wire \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/rx_tp_nump[3] ;
wire \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/rx_tp_nump[2] ;
wire \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/rx_tp_nump[1] ;
wire \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/rx_tp_nump[0] ;
wire \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/rx_tp_seq[4] ;
wire \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/rx_tp_seq[3] ;
wire \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/rx_tp_seq[2] ;
wire \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/rx_tp_seq[1] ;
wire \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/rx_tp_seq[0] ;
wire \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/rx_tp_stream[15] ;
wire \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/rx_tp_stream[14] ;
wire \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/rx_tp_stream[13] ;
wire \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/rx_tp_stream[12] ;
wire \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/rx_tp_stream[11] ;
wire \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/rx_tp_stream[10] ;
wire \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/rx_tp_stream[9] ;
wire \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/rx_tp_stream[8] ;
wire \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/rx_tp_stream[7] ;
wire \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/rx_tp_stream[6] ;
wire \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/rx_tp_stream[5] ;
wire \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/rx_tp_stream[4] ;
wire \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/rx_tp_stream[3] ;
wire \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/rx_tp_stream[2] ;
wire \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/rx_tp_stream[1] ;
wire \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/rx_tp_stream[0] ;
wire \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/rx_tp ;
wire \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/rx_tp_retry ;
wire \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/rx_tp_pktpend ;
wire \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/tx_tp_a_subtype[3] ;
wire \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/tx_tp_a_subtype[2] ;
wire \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/tx_tp_a_subtype[1] ;
wire \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/tx_tp_a_subtype[0] ;
wire \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/tx_tp_a_endp[3] ;
wire \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/tx_tp_a_endp[2] ;
wire \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/tx_tp_a_endp[1] ;
wire \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/tx_tp_a_endp[0] ;
wire \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/tx_tp_a ;
wire \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/tx_tp_a_dir ;
wire \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/tx_tp_a_nump[4] ;
wire \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/tx_tp_a_nump[3] ;
wire \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/tx_tp_a_nump[2] ;
wire \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/tx_tp_a_nump[1] ;
wire \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/tx_tp_a_nump[0] ;
wire \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/tx_tp_a_seq[4] ;
wire \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/tx_tp_a_seq[3] ;
wire \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/tx_tp_a_seq[2] ;
wire \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/tx_tp_a_seq[1] ;
wire \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/tx_tp_a_seq[0] ;
wire \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/tx_tp_a_stream[15] ;
wire \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/tx_tp_a_stream[14] ;
wire \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/tx_tp_a_stream[13] ;
wire \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/tx_tp_a_stream[12] ;
wire \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/tx_tp_a_stream[11] ;
wire \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/tx_tp_a_stream[10] ;
wire \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/tx_tp_a_stream[9] ;
wire \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/tx_tp_a_stream[8] ;
wire \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/tx_tp_a_stream[7] ;
wire \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/tx_tp_a_stream[6] ;
wire \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/tx_tp_a_stream[5] ;
wire \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/tx_tp_a_stream[4] ;
wire \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/tx_tp_a_stream[3] ;
wire \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/tx_tp_a_stream[2] ;
wire \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/tx_tp_a_stream[1] ;
wire \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/tx_tp_a_stream[0] ;
wire \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/tx_tp_a_retry ;
wire \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/tx_tp_b_subtype[3] ;
wire \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/tx_tp_b_subtype[2] ;
wire \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/tx_tp_b_subtype[1] ;
wire \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/tx_tp_b_subtype[0] ;
wire \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/tx_tp_b_endp[3] ;
wire \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/tx_tp_b_endp[2] ;
wire \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/tx_tp_b_endp[1] ;
wire \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/tx_tp_b_endp[0] ;
wire \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/tx_tp_b ;
wire \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/tx_tp_b_retry ;
wire \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/tx_tp_b_nump[4] ;
wire \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/tx_tp_b_nump[3] ;
wire \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/tx_tp_b_nump[2] ;
wire \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/tx_tp_b_nump[1] ;
wire \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/tx_tp_b_nump[0] ;
wire \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/tx_tp_c_subtype[3] ;
wire \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/tx_tp_c_subtype[2] ;
wire \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/tx_tp_c_subtype[1] ;
wire \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/tx_tp_c_subtype[0] ;
wire \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/tx_tp_c_endp[3] ;
wire \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/tx_tp_c_endp[2] ;
wire \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/tx_tp_c_endp[1] ;
wire \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/tx_tp_c_endp[0] ;
wire \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/tx_tp_c ;
wire \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/tx_tp_c_retry ;
wire \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/tx_tp_c_nump[4] ;
wire \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/tx_tp_c_nump[3] ;
wire \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/tx_tp_c_nump[2] ;
wire \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/tx_tp_c_nump[1] ;
wire \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/tx_tp_c_nump[0] ;
wire \UserLayer_top_inst/DataTransfer_inst/ep1_in_buf_ready ;
wire \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/iu3ep0/req_cnt[7] ;
wire \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/iu3ep0/req_cnt[6] ;
wire \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/iu3ep0/req_cnt[5] ;
wire \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/iu3ep0/req_cnt[4] ;
wire \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/iu3ep0/req_cnt[3] ;
wire \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/iu3ep0/req_cnt[2] ;
wire \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/iu3ep0/req_cnt[1] ;
wire \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/iu3ep0/req_cnt[0] ;
wire \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/host_requests_data ;
wire \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/host_requests_endpt[3] ;
wire \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/host_requests_endpt[2] ;
wire \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/host_requests_endpt[1] ;
wire \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/host_requests_endpt[0] ;
wire \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/rx_dpp_start ;
wire \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/rx_dpp_done ;
wire \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/rx_dpp_crcgood ;
wire \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/err_missed_dpp_start ;
wire \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/err_missed_dpp_done ;
wire \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/tx_dph ;
wire \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/tx_dph_eob ;
wire \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/tx_dph_dir ;
wire \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/tx_dph_endp[3] ;
wire \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/tx_dph_endp[2] ;
wire \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/tx_dph_endp[1] ;
wire \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/tx_dph_endp[0] ;
wire \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/tx_dph_seq[4] ;
wire \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/tx_dph_seq[3] ;
wire \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/tx_dph_seq[2] ;
wire \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/tx_dph_seq[1] ;
wire \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/tx_dph_seq[0] ;
wire \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/tx_dph_len[15] ;
wire \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/tx_dph_len[14] ;
wire \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/tx_dph_len[13] ;
wire \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/tx_dph_len[12] ;
wire \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/tx_dph_len[11] ;
wire \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/tx_dph_len[10] ;
wire \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/tx_dph_len[9] ;
wire \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/tx_dph_len[8] ;
wire \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/tx_dph_len[7] ;
wire \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/tx_dph_len[6] ;
wire \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/tx_dph_len[5] ;
wire \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/tx_dph_len[4] ;
wire \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/tx_dph_len[3] ;
wire \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/tx_dph_len[2] ;
wire \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/tx_dph_len[1] ;
wire \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/tx_dph_len[0] ;
wire \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/tx_dpp_ack ;
wire \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/tx_dpp_done ;
wire \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/ep2_buf_out_nump[4] ;
wire \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/ep2_buf_out_nump[3] ;
wire \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/ep2_buf_out_nump[2] ;
wire \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/ep2_buf_out_nump[1] ;
wire \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/ep2_buf_out_nump[0] ;
wire \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/burst_in_act ;
wire \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/burst_in_stop ;
wire \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/do_send_dpp ;
wire \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/do_send_dpp_ack ;
wire \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/do_send_dpp_eob ;
wire \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/crc_hprx_out[15] ;
wire \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/crc_hprx_out[14] ;
wire \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/crc_hprx_out[13] ;
wire \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/crc_hprx_out[12] ;
wire \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/crc_hprx_out[11] ;
wire \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/crc_hprx_out[10] ;
wire \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/crc_hprx_out[9] ;
wire \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/crc_hprx_out[8] ;
wire \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/crc_hprx_out[7] ;
wire \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/crc_hprx_out[6] ;
wire \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/crc_hprx_out[5] ;
wire \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/crc_hprx_out[4] ;
wire \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/crc_hprx_out[3] ;
wire \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/crc_hprx_out[2] ;
wire \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/crc_hprx_out[1] ;
wire \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/crc_hprx_out[0] ;
wire \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/crc_hprx_rst ;
wire \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/crc_hprx_en ;
wire \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/crc_hprx_in[31] ;
wire \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/crc_hprx_in[30] ;
wire \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/crc_hprx_in[29] ;
wire \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/crc_hprx_in[28] ;
wire \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/crc_hprx_in[27] ;
wire \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/crc_hprx_in[26] ;
wire \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/crc_hprx_in[25] ;
wire \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/crc_hprx_in[24] ;
wire \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/crc_hprx_in[23] ;
wire \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/crc_hprx_in[22] ;
wire \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/crc_hprx_in[21] ;
wire \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/crc_hprx_in[20] ;
wire \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/crc_hprx_in[19] ;
wire \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/crc_hprx_in[18] ;
wire \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/crc_hprx_in[17] ;
wire \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/crc_hprx_in[16] ;
wire \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/crc_hprx_in[15] ;
wire \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/crc_hprx_in[14] ;
wire \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/crc_hprx_in[13] ;
wire \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/crc_hprx_in[12] ;
wire \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/crc_hprx_in[11] ;
wire \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/crc_hprx_in[10] ;
wire \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/crc_hprx_in[9] ;
wire \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/crc_hprx_in[8] ;
wire \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/crc_hprx_in[7] ;
wire \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/crc_hprx_in[6] ;
wire \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/crc_hprx_in[5] ;
wire \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/crc_hprx_in[4] ;
wire \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/crc_hprx_in[3] ;
wire \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/crc_hprx_in[2] ;
wire \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/crc_hprx_in[1] ;
wire \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/crc_hprx_in[0] ;
wire \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/crc_cw3_out[4] ;
wire \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/crc_cw3_out[3] ;
wire \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/crc_cw3_out[2] ;
wire \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/crc_cw3_out[1] ;
wire \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/crc_cw3_out[0] ;
wire \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/in_header_cw[15] ;
wire \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/in_header_cw[14] ;
wire \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/in_header_cw[13] ;
wire \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/in_header_cw[12] ;
wire \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/in_header_cw[11] ;
wire \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/in_header_cw[10] ;
wire \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/in_header_cw[9] ;
wire \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/in_header_cw[8] ;
wire \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/in_header_cw[7] ;
wire \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/in_header_cw[6] ;
wire \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/in_header_cw[5] ;
wire \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/in_header_cw[4] ;
wire \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/in_header_cw[3] ;
wire \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/in_header_cw[2] ;
wire \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/in_header_cw[1] ;
wire \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/in_header_cw[0] ;
wire \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/in_link_command[10] ;
wire \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/in_link_command[9] ;
wire \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/in_link_command[8] ;
wire \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/in_link_command[7] ;
wire \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/in_link_command[6] ;
wire \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/in_link_command[5] ;
wire \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/in_link_command[4] ;
wire \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/in_link_command[3] ;
wire \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/in_link_command[2] ;
wire \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/in_link_command[1] ;
wire \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/in_link_command[0] ;
wire \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/crc_cw1_out[4] ;
wire \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/crc_cw1_out[3] ;
wire \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/crc_cw1_out[2] ;
wire \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/crc_cw1_out[1] ;
wire \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/crc_cw1_out[0] ;
wire \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/in_link_command[31] ;
wire \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/in_link_command[30] ;
wire \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/in_link_command[29] ;
wire \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/in_link_command[28] ;
wire \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/in_link_command[27] ;
wire \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/in_link_command[26] ;
wire \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/in_link_command[25] ;
wire \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/in_link_command[24] ;
wire \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/in_link_command[23] ;
wire \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/in_link_command[22] ;
wire \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/in_link_command[21] ;
wire \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/in_link_command[20] ;
wire \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/in_link_command[19] ;
wire \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/in_link_command[18] ;
wire \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/in_link_command[17] ;
wire \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/in_link_command[16] ;
wire \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/crc_cw2_out[4] ;
wire \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/crc_cw2_out[3] ;
wire \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/crc_cw2_out[2] ;
wire \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/crc_cw2_out[1] ;
wire \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/crc_cw2_out[0] ;
wire \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/in_link_command[15] ;
wire \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/in_link_command[14] ;
wire \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/in_link_command[13] ;
wire \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/in_link_command[12] ;
wire \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/in_link_command[11] ;
wire \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/err_lbad_reg ;
wire \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/rx_hdr_seq_num_reg[2] ;
wire \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/rx_hdr_seq_num_reg[1] ;
wire \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/rx_hdr_seq_num_reg[0] ;
wire \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/link_err ;
wire \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/tx_lbad_pop ;
wire \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/tx_lbad_q[10] ;
wire \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/tx_lbad_q[9] ;
wire \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/tx_lbad_q[8] ;
wire \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/tx_lbad_q[7] ;
wire \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/tx_lbad_q[6] ;
wire \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/tx_lbad_q[5] ;
wire \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/tx_lbad_q[4] ;
wire \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/tx_lbad_q[3] ;
wire \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/tx_lbad_q[2] ;
wire \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/tx_lbad_q[1] ;
wire \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/tx_lbad_q[0] ;
wire \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/tx_lbad_empty ;
wire \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/tx_lbad_act ;
wire \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/wait_retry ;
wire \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/rx_retry ;
wire \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/hp_valid_k_cnt[2] ;
wire \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/hp_valid_k_cnt[1] ;
wire \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/hp_valid_k_cnt[0] ;
wire \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/hp_valid_k[3] ;
wire \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/hp_valid_k[2] ;
wire \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/hp_valid_k[1] ;
wire \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/hp_valid_k[0] ;
wire \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/queue_state[2] ;
wire \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/queue_state[1] ;
wire \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/queue_state[0] ;
wire \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/send_dpp_state[3] ;
wire \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/send_dpp_state[2] ;
wire \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/send_dpp_state[1] ;
wire \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/send_dpp_state[0] ;
wire \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/tx_link_busy ;
wire \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/tx_lcmd_req ;
wire \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/tx_hp_req ;
wire \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/ltssm_state[4] ;
wire \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/ltssm_state[3] ;
wire \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/ltssm_state[2] ;
wire \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/ltssm_state[1] ;
wire \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/ltssm_state[0] ;
wire \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/reset_n ;
wire \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/ltssm_go_recovery ;
wire \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/res_mem_wr_en ;
wire \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/res_mem_wr_dat[35] ;
wire \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/res_mem_wr_dat[34] ;
wire \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/res_mem_wr_dat[33] ;
wire \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/res_mem_wr_dat[32] ;
wire \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/res_mem_wr_dat[31] ;
wire \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/res_mem_wr_dat[30] ;
wire \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/res_mem_wr_dat[29] ;
wire \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/res_mem_wr_dat[28] ;
wire \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/res_mem_wr_dat[27] ;
wire \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/res_mem_wr_dat[26] ;
wire \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/res_mem_wr_dat[25] ;
wire \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/res_mem_wr_dat[24] ;
wire \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/res_mem_wr_dat[23] ;
wire \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/res_mem_wr_dat[22] ;
wire \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/res_mem_wr_dat[21] ;
wire \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/res_mem_wr_dat[20] ;
wire \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/res_mem_wr_dat[19] ;
wire \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/res_mem_wr_dat[18] ;
wire \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/res_mem_wr_dat[17] ;
wire \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/res_mem_wr_dat[16] ;
wire \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/res_mem_wr_dat[15] ;
wire \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/res_mem_wr_dat[14] ;
wire \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/res_mem_wr_dat[13] ;
wire \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/res_mem_wr_dat[12] ;
wire \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/res_mem_wr_dat[11] ;
wire \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/res_mem_wr_dat[10] ;
wire \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/res_mem_wr_dat[9] ;
wire \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/res_mem_wr_dat[8] ;
wire \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/res_mem_wr_dat[7] ;
wire \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/res_mem_wr_dat[6] ;
wire \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/res_mem_wr_dat[5] ;
wire \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/res_mem_wr_dat[4] ;
wire \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/res_mem_wr_dat[3] ;
wire \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/res_mem_wr_dat[2] ;
wire \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/res_mem_wr_dat[1] ;
wire \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/res_mem_wr_dat[0] ;
wire \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/res_mem_wr_addr[10] ;
wire \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/res_mem_wr_addr[9] ;
wire \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/res_mem_wr_addr[8] ;
wire \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/res_mem_wr_addr[7] ;
wire \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/res_mem_wr_addr[6] ;
wire \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/res_mem_wr_addr[5] ;
wire \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/res_mem_wr_addr[4] ;
wire \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/res_mem_wr_addr[3] ;
wire \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/res_mem_wr_addr[2] ;
wire \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/res_mem_wr_addr[1] ;
wire \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/res_mem_wr_addr[0] ;
wire \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/res_mem_wr_pt[1] ;
wire \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/res_mem_wr_pt[0] ;
wire \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/resend_hp_act ;
wire \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/tx_hdr_seq_num_dec[2] ;
wire \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/tx_hdr_seq_num_dec[1] ;
wire \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/tx_hdr_seq_num_dec[0] ;
wire \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/resend_hp_num[4] ;
wire \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/resend_hp_num[3] ;
wire \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/resend_hp_num[2] ;
wire \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/resend_hp_num[1] ;
wire \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/resend_hp_num[0] ;
wire \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/res_mem_rd_pt[1] ;
wire \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/res_mem_rd_pt[0] ;
wire \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/res_mem_rd_addr[10] ;
wire \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/res_mem_rd_addr[9] ;
wire \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/res_mem_rd_addr[8] ;
wire \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/res_mem_rd_addr[7] ;
wire \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/res_mem_rd_addr[6] ;
wire \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/res_mem_rd_addr[5] ;
wire \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/res_mem_rd_addr[4] ;
wire \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/res_mem_rd_addr[3] ;
wire \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/res_mem_rd_addr[2] ;
wire \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/res_mem_rd_addr[1] ;
wire \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/res_mem_rd_addr[0] ;
wire \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/res_mem_rd_en ;
wire \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/tx_res_req ;
wire \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/tx_res_req_ack ;
wire \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/res_mem_rd_dat[35] ;
wire \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/res_mem_rd_dat[34] ;
wire \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/res_mem_rd_dat[33] ;
wire \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/res_mem_rd_dat[32] ;
wire \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/res_mem_rd_dat[31] ;
wire \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/res_mem_rd_dat[30] ;
wire \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/res_mem_rd_dat[29] ;
wire \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/res_mem_rd_dat[28] ;
wire \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/res_mem_rd_dat[27] ;
wire \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/res_mem_rd_dat[26] ;
wire \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/res_mem_rd_dat[25] ;
wire \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/res_mem_rd_dat[24] ;
wire \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/res_mem_rd_dat[23] ;
wire \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/res_mem_rd_dat[22] ;
wire \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/res_mem_rd_dat[21] ;
wire \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/res_mem_rd_dat[20] ;
wire \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/res_mem_rd_dat[19] ;
wire \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/res_mem_rd_dat[18] ;
wire \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/res_mem_rd_dat[17] ;
wire \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/res_mem_rd_dat[16] ;
wire \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/res_mem_rd_dat[15] ;
wire \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/res_mem_rd_dat[14] ;
wire \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/res_mem_rd_dat[13] ;
wire \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/res_mem_rd_dat[12] ;
wire \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/res_mem_rd_dat[11] ;
wire \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/res_mem_rd_dat[10] ;
wire \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/res_mem_rd_dat[9] ;
wire \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/res_mem_rd_dat[8] ;
wire \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/res_mem_rd_dat[7] ;
wire \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/res_mem_rd_dat[6] ;
wire \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/res_mem_rd_dat[5] ;
wire \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/res_mem_rd_dat[4] ;
wire \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/res_mem_rd_dat[3] ;
wire \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/res_mem_rd_dat[2] ;
wire \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/res_mem_rd_dat[1] ;
wire \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/res_mem_rd_dat[0] ;
wire \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/res_mem_rd_dat_val ;
wire \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/out_data_5[31] ;
wire \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/out_data_5[30] ;
wire \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/out_data_5[29] ;
wire \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/out_data_5[28] ;
wire \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/out_data_5[27] ;
wire \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/out_data_5[26] ;
wire \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/out_data_5[25] ;
wire \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/out_data_5[24] ;
wire \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/out_data_5[23] ;
wire \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/out_data_5[22] ;
wire \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/out_data_5[21] ;
wire \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/out_data_5[20] ;
wire \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/out_data_5[19] ;
wire \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/out_data_5[18] ;
wire \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/out_data_5[17] ;
wire \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/out_data_5[16] ;
wire \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/out_data_5[15] ;
wire \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/out_data_5[14] ;
wire \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/out_data_5[13] ;
wire \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/out_data_5[12] ;
wire \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/out_data_5[11] ;
wire \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/out_data_5[10] ;
wire \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/out_data_5[9] ;
wire \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/out_data_5[8] ;
wire \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/out_data_5[7] ;
wire \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/out_data_5[6] ;
wire \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/out_data_5[5] ;
wire \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/out_data_5[4] ;
wire \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/out_data_5[3] ;
wire \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/out_data_5[2] ;
wire \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/out_data_5[1] ;
wire \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/out_data_5[0] ;
wire \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/out_datak_5[3] ;
wire \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/out_datak_5[2] ;
wire \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/out_datak_5[1] ;
wire \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/out_datak_5[0] ;
wire \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/out_active_5 ;
wire \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/tx_hdr_seq_num_dec_latch[2] ;
wire \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/tx_hdr_seq_num_dec_latch[1] ;
wire \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/tx_hdr_seq_num_dec_latch[0] ;
wire \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/tx_lgood_empty ;
wire \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/tx_lcrd_empty ;
wire \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/send_hp_state[2] ;
wire \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/send_hp_state[1] ;
wire \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/send_hp_state[0] ;
wire \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/send_lcmd_state[3] ;
wire \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/send_lcmd_state[2] ;
wire \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/send_lcmd_state[1] ;
wire \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/send_lcmd_state[0] ;
wire \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/tx_sel[2] ;
wire \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/tx_sel[1] ;
wire \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/tx_sel[0] ;
wire \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/tx_lcrd_act ;
wire \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/qc[7] ;
wire \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/qc[6] ;
wire \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/qc[5] ;
wire \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/qc[4] ;
wire \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/qc[3] ;
wire \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/qc[2] ;
wire \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/qc[1] ;
wire \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/qc[0] ;
wire \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/tx_lgood_act ;
wire \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/res_state[2] ;
wire \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/res_state[1] ;
wire \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/res_state[0] ;
wire \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/buf_out_dp_acked[2] ;
wire \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/usb3_ep2_IN/buf_in_ready ;
wire \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/usb3_ep2_IN/buf_in_commit ;
wire \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/usb3_ep2_IN/buf_in_eob ;
wire \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/usb3_ep2_IN/in_ep_rty ;
wire \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/usb3_ep2_IN/buf_out_hasdata ;
wire \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/usb3_ep2_IN/buf_out_eob ;
wire \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/usb3_ep2_IN/buf_out_nump[4] ;
wire \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/usb3_ep2_IN/buf_out_nump[3] ;
wire \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/usb3_ep2_IN/buf_out_nump[2] ;
wire \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/usb3_ep2_IN/buf_out_nump[1] ;
wire \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/usb3_ep2_IN/buf_out_nump[0] ;
wire \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/usb3_ep2_IN/buf_out_next_dp_ack_pt[3] ;
wire \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/usb3_ep2_IN/buf_out_next_dp_ack_pt[2] ;
wire \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/usb3_ep2_IN/buf_out_next_dp_ack_pt[1] ;
wire \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/usb3_ep2_IN/buf_out_next_dp_ack_pt[0] ;
wire \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/usb3_ep2_IN/buf_wt_ack_mem[15] ;
wire \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/usb3_ep2_IN/buf_wt_ack_mem[14] ;
wire \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/usb3_ep2_IN/buf_wt_ack_mem[13] ;
wire \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/usb3_ep2_IN/buf_wt_ack_mem[12] ;
wire \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/usb3_ep2_IN/buf_wt_ack_mem[11] ;
wire \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/usb3_ep2_IN/buf_wt_ack_mem[10] ;
wire \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/usb3_ep2_IN/buf_wt_ack_mem[9] ;
wire \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/usb3_ep2_IN/buf_wt_ack_mem[8] ;
wire \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/usb3_ep2_IN/buf_wt_ack_mem[7] ;
wire \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/usb3_ep2_IN/buf_wt_ack_mem[6] ;
wire \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/usb3_ep2_IN/buf_wt_ack_mem[5] ;
wire \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/usb3_ep2_IN/buf_wt_ack_mem[4] ;
wire \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/usb3_ep2_IN/buf_wt_ack_mem[3] ;
wire \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/usb3_ep2_IN/buf_wt_ack_mem[2] ;
wire \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/usb3_ep2_IN/buf_wt_ack_mem[1] ;
wire \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/usb3_ep2_IN/buf_wt_ack_mem[0] ;
wire \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/usb3_ep2_IN/buf_ready_mem[0] ;
wire \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/usb3_ep2_IN/buf_ready_mem[1] ;
wire \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/usb3_ep2_IN/buf_ready_mem[2] ;
wire \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/usb3_ep2_IN/buf_ready_mem[3] ;
wire \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/usb3_ep2_IN/buf_ready_mem[4] ;
wire \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/usb3_ep2_IN/buf_ready_mem[5] ;
wire \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/usb3_ep2_IN/buf_ready_mem[6] ;
wire \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/usb3_ep2_IN/buf_ready_mem[7] ;
wire \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/usb3_ep2_IN/buf_ready_mem[8] ;
wire \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/usb3_ep2_IN/buf_ready_mem[9] ;
wire \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/usb3_ep2_IN/buf_ready_mem[10] ;
wire \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/usb3_ep2_IN/buf_ready_mem[11] ;
wire \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/usb3_ep2_IN/buf_ready_mem[12] ;
wire \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/usb3_ep2_IN/buf_ready_mem[13] ;
wire \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/usb3_ep2_IN/buf_ready_mem[14] ;
wire \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/usb3_ep2_IN/buf_ready_mem[15] ;
wire \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/usb3_ep2_IN/buf_out_hasdata_mem[0] ;
wire \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/usb3_ep2_IN/buf_out_hasdata_mem[1] ;
wire \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/usb3_ep2_IN/buf_out_hasdata_mem[2] ;
wire \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/usb3_ep2_IN/buf_out_hasdata_mem[3] ;
wire \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/usb3_ep2_IN/buf_out_hasdata_mem[4] ;
wire \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/usb3_ep2_IN/buf_out_hasdata_mem[5] ;
wire \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/usb3_ep2_IN/buf_out_hasdata_mem[6] ;
wire \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/usb3_ep2_IN/buf_out_hasdata_mem[7] ;
wire \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/usb3_ep2_IN/buf_out_hasdata_mem[8] ;
wire \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/usb3_ep2_IN/buf_out_hasdata_mem[9] ;
wire \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/usb3_ep2_IN/buf_out_hasdata_mem[10] ;
wire \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/usb3_ep2_IN/buf_out_hasdata_mem[11] ;
wire \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/usb3_ep2_IN/buf_out_hasdata_mem[12] ;
wire \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/usb3_ep2_IN/buf_out_hasdata_mem[13] ;
wire \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/usb3_ep2_IN/buf_out_hasdata_mem[14] ;
wire \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/usb3_ep2_IN/buf_out_hasdata_mem[15] ;
wire \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/err_lbad_recv_latch ;
wire \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/err_lbad_recv_latch_2 ;
wire \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/usb3_ep2_IN/buf_out_pt[3] ;
wire \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/usb3_ep2_IN/buf_out_pt[2] ;
wire \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/usb3_ep2_IN/buf_out_pt[1] ;
wire \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/usb3_ep2_IN/buf_out_pt[0] ;
wire \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/usb3_ep2_IN/buf_in_pt[3] ;
wire \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/usb3_ep2_IN/buf_in_pt[2] ;
wire \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/usb3_ep2_IN/buf_in_pt[1] ;
wire \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/usb3_ep2_IN/buf_in_pt[0] ;
wire \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/usb3_ep2_IN/wt_ack_pt[3] ;
wire \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/usb3_ep2_IN/wt_ack_pt[2] ;
wire \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/usb3_ep2_IN/wt_ack_pt[1] ;
wire \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/usb3_ep2_IN/wt_ack_pt[0] ;
wire \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/tx_hp_act ;
wire \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/err_hp_seq_latch ;
wire \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/err_lgood_order_latch ;
wire \USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/tx_lgood_pop ;
wire request_active;
wire ep2_in_buf_data_commit;
wire ep2_in_buf_eob;
wire \UserLayer_top_inst/cam_active ;
wire \dbg_ltssm_state[4] ;
wire \dbg_ltssm_state[3] ;
wire \dbg_ltssm_state[2] ;
wire \dbg_ltssm_state[1] ;
wire \dbg_ltssm_state[0] ;
wire pclk;
wire tms_pad_i;
wire tck_pad_i;
wire tdi_pad_i;
wire tdo_pad_o;
wire tms_i_c;
wire tck_i_c;
wire tdi_i_c;
wire tdo_o_c;
wire [9:0] control0;
wire gao_jtag_tck;
wire gao_jtag_reset;
wire run_test_idle_er1;
wire run_test_idle_er2;
wire shift_dr_capture_dr;
wire update_dr;
wire pause_dr;
wire enable_er1;
wire enable_er2;
wire gao_jtag_tdi;
wire tdo_er1;

IBUF tms_ibuf (
    .I(tms_pad_i),
    .O(tms_i_c)
);

IBUF tck_ibuf (
    .I(tck_pad_i),
    .O(tck_i_c)
);

IBUF tdi_ibuf (
    .I(tdi_pad_i),
    .O(tdi_i_c)
);

OBUF tdo_obuf (
    .I(tdo_o_c),
    .O(tdo_pad_o)
);

GW_JTAG  u_gw_jtag(
    .tms_pad_i(tms_i_c),
    .tck_pad_i(tck_i_c),
    .tdi_pad_i(tdi_i_c),
    .tdo_pad_o(tdo_o_c),
    .tck_o(gao_jtag_tck),
    .test_logic_reset_o(gao_jtag_reset),
    .run_test_idle_er1_o(run_test_idle_er1),
    .run_test_idle_er2_o(run_test_idle_er2),
    .shift_dr_capture_dr_o(shift_dr_capture_dr),
    .update_dr_o(update_dr),
    .pause_dr_o(pause_dr),
    .enable_er1_o(enable_er1),
    .enable_er2_o(enable_er2),
    .tdi_o(gao_jtag_tdi),
    .tdo_er1_i(tdo_er1),
    .tdo_er2_i(1'b0)
);

gw_con_top  u_icon_top(
    .tck_i(gao_jtag_tck),
    .tdi_i(gao_jtag_tdi),
    .tdo_o(tdo_er1),
    .rst_i(gao_jtag_reset),
    .control0(control0[9:0]),
    .enable_i(enable_er1),
    .shift_dr_capture_dr_i(shift_dr_capture_dr),
    .update_dr_i(update_dr)
);

ao_top_0  u_la0_top(
    .control(control0[9:0]),
    .trig0_i(request_active),
    .trig1_i({ep2_in_buf_data_commit,ep2_in_buf_eob}),
    .trig2_i({\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/host_requests_endpt[3] ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/host_requests_endpt[2] ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/host_requests_endpt[1] ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/host_requests_endpt[0] }),
    .trig3_i(\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/host_requests_data ),
    .trig4_i(\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/buf_out_dp_acked[2] ),
    .trig5_i({\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/tx_dph ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/tx_dph_eob }),
    .trig6_i(\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/rx_tp_retry ),
    .trig7_i({\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/rx_tp ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/rx_tp_endp[3] ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/rx_tp_endp[2] ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/rx_tp_endp[1] ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/rx_tp_endp[0] }),
    .trig8_i({\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/err_lbad_reg ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/link_err ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/burst_in_act ,\UserLayer_top_inst/cam_active ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/err_lgood_order ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/err_hp_seq ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/err_lbad_recv }),
    .trig9_i({\dbg_ltssm_state[4] ,\dbg_ltssm_state[3] ,\dbg_ltssm_state[2] ,\dbg_ltssm_state[1] ,\dbg_ltssm_state[0] }),
    .data_i({\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/in_data[31] ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/in_data[30] ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/in_data[29] ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/in_data[28] ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/in_data[27] ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/in_data[26] ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/in_data[25] ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/in_data[24] ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/in_data[23] ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/in_data[22] ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/in_data[21] ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/in_data[20] ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/in_data[19] ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/in_data[18] ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/in_data[17] ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/in_data[16] ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/in_data[15] ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/in_data[14] ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/in_data[13] ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/in_data[12] ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/in_data[11] ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/in_data[10] ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/in_data[9] ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/in_data[8] ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/in_data[7] ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/in_data[6] ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/in_data[5] ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/in_data[4] ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/in_data[3] ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/in_data[2] ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/in_data[1] ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/in_data[0] ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/in_datak[3] ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/in_datak[2] ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/in_datak[1] ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/in_datak[0] ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/in_active ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/outp_data[31] ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/outp_data[30] ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/outp_data[29] ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/outp_data[28] ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/outp_data[27] ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/outp_data[26] ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/outp_data[25] ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/outp_data[24] ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/outp_data[23] ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/outp_data[22] ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/outp_data[21] ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/outp_data[20] ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/outp_data[19] ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/outp_data[18] ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/outp_data[17] ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/outp_data[16] ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/outp_data[15] ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/outp_data[14] ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/outp_data[13] ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/outp_data[12] ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/outp_data[11] ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/outp_data[10] ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/outp_data[9] ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/outp_data[8] ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/outp_data[7] ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/outp_data[6] ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/outp_data[5] ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/outp_data[4] ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/outp_data[3] ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/outp_data[2] ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/outp_data[1] ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/outp_data[0] ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/outp_datak[3] ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/outp_datak[2] ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/outp_datak[1] ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/outp_datak[0] ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/outp_active ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/out_stall ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/enter_u0_cnt[7] ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/enter_u0_cnt[6] ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/enter_u0_cnt[5] ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/enter_u0_cnt[4] ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/enter_u0_cnt[3] ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/enter_u0_cnt[2] ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/enter_u0_cnt[1] ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/enter_u0_cnt[0] ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/ltssm_exit_u0 ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/ltssm_current_state[4] ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/ltssm_current_state[3] ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/ltssm_current_state[2] ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/ltssm_current_state[1] ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/ltssm_current_state[0] ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/queue_send_u0_adv ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/queue_send_u0_portcap ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/link_cmd_det ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/send_port_cfg_resp ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/remote_rx_cred_count[2] ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/remote_rx_cred_count[1] ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/remote_rx_cred_count[0] ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/tx_cred_idx[1] ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/tx_cred_idx[0] ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/send_port_cfg_resp_ack ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/ack_tx_hdr_seq_num[2] ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/ack_tx_hdr_seq_num[1] ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/ack_tx_hdr_seq_num[0] ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/rx_hdr_seq_num[2] ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/rx_hdr_seq_num[1] ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/rx_hdr_seq_num[0] ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/ltssm_enter_u0_by_polling ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/in_link_command_act ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/in_link_command_crc_good ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/in_link_command_latch_act ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/recv_u0_adv ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/err_lgood_order ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/err_lcrd_mismatch ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/err_lbad_recv ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/hp_det ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/in_header_act ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/hp_crc_good ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/err_hp_seq ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/err_lbad ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/local_rx_cred_count[2] ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/local_rx_cred_count[1] ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/local_rx_cred_count[0] ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/rx_dph ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/rx_dph_eob ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/rx_dph_setup ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/rx_dph_pktpend ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/rx_dph_endp[3] ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/rx_dph_endp[2] ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/rx_dph_endp[1] ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/rx_dph_endp[0] ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/rx_dph_seq[4] ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/rx_dph_seq[3] ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/rx_dph_seq[2] ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/rx_dph_seq[1] ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/rx_dph_seq[0] ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/rx_dph_len[15] ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/rx_dph_len[14] ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/rx_dph_len[13] ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/rx_dph_len[12] ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/rx_dph_len[11] ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/rx_dph_len[10] ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/rx_dph_len[9] ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/rx_dph_len[8] ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/rx_dph_len[7] ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/rx_dph_len[6] ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/rx_dph_len[5] ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/rx_dph_len[4] ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/rx_dph_len[3] ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/rx_dph_len[2] ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/rx_dph_len[1] ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/rx_dph_len[0] ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/rx_tp_subtype[3] ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/rx_tp_subtype[2] ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/rx_tp_subtype[1] ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/rx_tp_subtype[0] ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/rx_tp_endp[3] ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/rx_tp_endp[2] ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/rx_tp_endp[1] ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/rx_tp_endp[0] ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/rx_tp_nump[4] ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/rx_tp_nump[3] ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/rx_tp_nump[2] ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/rx_tp_nump[1] ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/rx_tp_nump[0] ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/rx_tp_seq[4] ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/rx_tp_seq[3] ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/rx_tp_seq[2] ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/rx_tp_seq[1] ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/rx_tp_seq[0] ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/rx_tp_stream[15] ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/rx_tp_stream[14] ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/rx_tp_stream[13] ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/rx_tp_stream[12] ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/rx_tp_stream[11] ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/rx_tp_stream[10] ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/rx_tp_stream[9] ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/rx_tp_stream[8] ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/rx_tp_stream[7] ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/rx_tp_stream[6] ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/rx_tp_stream[5] ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/rx_tp_stream[4] ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/rx_tp_stream[3] ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/rx_tp_stream[2] ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/rx_tp_stream[1] ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/rx_tp_stream[0] ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/rx_tp ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/rx_tp_retry ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/rx_tp_pktpend ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/tx_tp_a_subtype[3] ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/tx_tp_a_subtype[2] ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/tx_tp_a_subtype[1] ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/tx_tp_a_subtype[0] ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/tx_tp_a_endp[3] ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/tx_tp_a_endp[2] ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/tx_tp_a_endp[1] ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/tx_tp_a_endp[0] ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/tx_tp_a ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/tx_tp_a_dir ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/tx_tp_a_nump[4] ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/tx_tp_a_nump[3] ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/tx_tp_a_nump[2] ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/tx_tp_a_nump[1] ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/tx_tp_a_nump[0] ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/tx_tp_a_seq[4] ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/tx_tp_a_seq[3] ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/tx_tp_a_seq[2] ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/tx_tp_a_seq[1] ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/tx_tp_a_seq[0] ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/tx_tp_a_stream[15] ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/tx_tp_a_stream[14] ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/tx_tp_a_stream[13] ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/tx_tp_a_stream[12] ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/tx_tp_a_stream[11] ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/tx_tp_a_stream[10] ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/tx_tp_a_stream[9] ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/tx_tp_a_stream[8] ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/tx_tp_a_stream[7] ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/tx_tp_a_stream[6] ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/tx_tp_a_stream[5] ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/tx_tp_a_stream[4] ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/tx_tp_a_stream[3] ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/tx_tp_a_stream[2] ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/tx_tp_a_stream[1] ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/tx_tp_a_stream[0] ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/tx_tp_a_retry ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/tx_tp_b_subtype[3] ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/tx_tp_b_subtype[2] ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/tx_tp_b_subtype[1] ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/tx_tp_b_subtype[0] ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/tx_tp_b_endp[3] ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/tx_tp_b_endp[2] ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/tx_tp_b_endp[1] ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/tx_tp_b_endp[0] ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/tx_tp_b ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/tx_tp_b_retry ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/tx_tp_b_nump[4] ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/tx_tp_b_nump[3] ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/tx_tp_b_nump[2] ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/tx_tp_b_nump[1] ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/tx_tp_b_nump[0] ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/tx_tp_c_subtype[3] ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/tx_tp_c_subtype[2] ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/tx_tp_c_subtype[1] ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/tx_tp_c_subtype[0] ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/tx_tp_c_endp[3] ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/tx_tp_c_endp[2] ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/tx_tp_c_endp[1] ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/tx_tp_c_endp[0] ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/tx_tp_c ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/tx_tp_c_retry ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/tx_tp_c_nump[4] ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/tx_tp_c_nump[3] ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/tx_tp_c_nump[2] ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/tx_tp_c_nump[1] ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/tx_tp_c_nump[0] ,\UserLayer_top_inst/DataTransfer_inst/ep1_in_buf_ready ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/iu3ep0/req_cnt[7] ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/iu3ep0/req_cnt[6] ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/iu3ep0/req_cnt[5] ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/iu3ep0/req_cnt[4] ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/iu3ep0/req_cnt[3] ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/iu3ep0/req_cnt[2] ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/iu3ep0/req_cnt[1] ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/iu3ep0/req_cnt[0] ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/host_requests_data ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/host_requests_endpt[3] ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/host_requests_endpt[2] ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/host_requests_endpt[1] ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/host_requests_endpt[0] ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/rx_dpp_start ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/rx_dpp_done ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/rx_dpp_crcgood ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/err_missed_dpp_start ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/err_missed_dpp_done ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/tx_dph ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/tx_dph_eob ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/tx_dph_dir ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/tx_dph_endp[3] ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/tx_dph_endp[2] ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/tx_dph_endp[1] ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/tx_dph_endp[0] ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/tx_dph_seq[4] ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/tx_dph_seq[3] ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/tx_dph_seq[2] ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/tx_dph_seq[1] ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/tx_dph_seq[0] ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/tx_dph_len[15] ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/tx_dph_len[14] ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/tx_dph_len[13] ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/tx_dph_len[12] ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/tx_dph_len[11] ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/tx_dph_len[10] ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/tx_dph_len[9] ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/tx_dph_len[8] ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/tx_dph_len[7] ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/tx_dph_len[6] ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/tx_dph_len[5] ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/tx_dph_len[4] ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/tx_dph_len[3] ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/tx_dph_len[2] ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/tx_dph_len[1] ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/tx_dph_len[0] ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/tx_dpp_ack ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/tx_dpp_done ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/ep2_buf_out_nump[4] ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/ep2_buf_out_nump[3] ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/ep2_buf_out_nump[2] ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/ep2_buf_out_nump[1] ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/ep2_buf_out_nump[0] ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/burst_in_act ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/burst_in_stop ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/do_send_dpp ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/do_send_dpp_ack ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/do_send_dpp_eob ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/crc_hprx_out[15] ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/crc_hprx_out[14] ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/crc_hprx_out[13] ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/crc_hprx_out[12] ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/crc_hprx_out[11] ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/crc_hprx_out[10] ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/crc_hprx_out[9] ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/crc_hprx_out[8] ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/crc_hprx_out[7] ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/crc_hprx_out[6] ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/crc_hprx_out[5] ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/crc_hprx_out[4] ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/crc_hprx_out[3] ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/crc_hprx_out[2] ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/crc_hprx_out[1] ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/crc_hprx_out[0] ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/crc_hprx_rst ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/crc_hprx_en ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/crc_hprx_in[31] ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/crc_hprx_in[30] ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/crc_hprx_in[29] ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/crc_hprx_in[28] ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/crc_hprx_in[27] ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/crc_hprx_in[26] ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/crc_hprx_in[25] ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/crc_hprx_in[24] ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/crc_hprx_in[23] ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/crc_hprx_in[22] ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/crc_hprx_in[21] ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/crc_hprx_in[20] ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/crc_hprx_in[19] ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/crc_hprx_in[18] ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/crc_hprx_in[17] ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/crc_hprx_in[16] ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/crc_hprx_in[15] ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/crc_hprx_in[14] ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/crc_hprx_in[13] ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/crc_hprx_in[12] ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/crc_hprx_in[11] ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/crc_hprx_in[10] ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/crc_hprx_in[9] ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/crc_hprx_in[8] ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/crc_hprx_in[7] ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/crc_hprx_in[6] ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/crc_hprx_in[5] ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/crc_hprx_in[4] ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/crc_hprx_in[3] ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/crc_hprx_in[2] ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/crc_hprx_in[1] ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/crc_hprx_in[0] ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/crc_cw3_out[4] ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/crc_cw3_out[3] ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/crc_cw3_out[2] ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/crc_cw3_out[1] ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/crc_cw3_out[0] ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/in_header_cw[15] ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/in_header_cw[14] ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/in_header_cw[13] ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/in_header_cw[12] ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/in_header_cw[11] ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/in_header_cw[10] ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/in_header_cw[9] ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/in_header_cw[8] ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/in_header_cw[7] ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/in_header_cw[6] ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/in_header_cw[5] ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/in_header_cw[4] ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/in_header_cw[3] ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/in_header_cw[2] ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/in_header_cw[1] ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/in_header_cw[0] ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/in_link_command[10] ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/in_link_command[9] ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/in_link_command[8] ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/in_link_command[7] ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/in_link_command[6] ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/in_link_command[5] ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/in_link_command[4] ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/in_link_command[3] ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/in_link_command[2] ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/in_link_command[1] ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/in_link_command[0] ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/crc_cw1_out[4] ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/crc_cw1_out[3] ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/crc_cw1_out[2] ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/crc_cw1_out[1] ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/crc_cw1_out[0] ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/in_link_command[31] ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/in_link_command[30] ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/in_link_command[29] ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/in_link_command[28] ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/in_link_command[27] ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/in_link_command[26] ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/in_link_command[25] ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/in_link_command[24] ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/in_link_command[23] ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/in_link_command[22] ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/in_link_command[21] ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/in_link_command[20] ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/in_link_command[19] ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/in_link_command[18] ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/in_link_command[17] ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/in_link_command[16] ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/crc_cw2_out[4] ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/crc_cw2_out[3] ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/crc_cw2_out[2] ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/crc_cw2_out[1] ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/crc_cw2_out[0] ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/in_link_command[15] ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/in_link_command[14] ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/in_link_command[13] ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/in_link_command[12] ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/in_link_command[11] ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/err_lbad_reg ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/rx_hdr_seq_num_reg[2] ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/rx_hdr_seq_num_reg[1] ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/rx_hdr_seq_num_reg[0] ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/link_err ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/tx_lbad_pop ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/tx_lbad_q[10] ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/tx_lbad_q[9] ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/tx_lbad_q[8] ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/tx_lbad_q[7] ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/tx_lbad_q[6] ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/tx_lbad_q[5] ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/tx_lbad_q[4] ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/tx_lbad_q[3] ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/tx_lbad_q[2] ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/tx_lbad_q[1] ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/tx_lbad_q[0] ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/tx_lbad_empty ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/tx_lbad_act ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/wait_retry ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/rx_retry ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/hp_valid_k_cnt[2] ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/hp_valid_k_cnt[1] ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/hp_valid_k_cnt[0] ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/hp_valid_k[3] ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/hp_valid_k[2] ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/hp_valid_k[1] ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/hp_valid_k[0] ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/queue_state[2] ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/queue_state[1] ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/queue_state[0] ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/send_dpp_state[3] ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/send_dpp_state[2] ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/send_dpp_state[1] ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/send_dpp_state[0] ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/tx_link_busy ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/tx_lcmd_req ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/tx_hp_req ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/ltssm_state[4] ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/ltssm_state[3] ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/ltssm_state[2] ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/ltssm_state[1] ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/ltssm_state[0] ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/reset_n ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/ltssm_go_recovery ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/res_mem_wr_en ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/res_mem_wr_dat[35] ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/res_mem_wr_dat[34] ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/res_mem_wr_dat[33] ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/res_mem_wr_dat[32] ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/res_mem_wr_dat[31] ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/res_mem_wr_dat[30] ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/res_mem_wr_dat[29] ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/res_mem_wr_dat[28] ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/res_mem_wr_dat[27] ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/res_mem_wr_dat[26] ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/res_mem_wr_dat[25] ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/res_mem_wr_dat[24] ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/res_mem_wr_dat[23] ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/res_mem_wr_dat[22] ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/res_mem_wr_dat[21] ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/res_mem_wr_dat[20] ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/res_mem_wr_dat[19] ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/res_mem_wr_dat[18] ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/res_mem_wr_dat[17] ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/res_mem_wr_dat[16] ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/res_mem_wr_dat[15] ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/res_mem_wr_dat[14] ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/res_mem_wr_dat[13] ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/res_mem_wr_dat[12] ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/res_mem_wr_dat[11] ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/res_mem_wr_dat[10] ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/res_mem_wr_dat[9] ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/res_mem_wr_dat[8] ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/res_mem_wr_dat[7] ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/res_mem_wr_dat[6] ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/res_mem_wr_dat[5] ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/res_mem_wr_dat[4] ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/res_mem_wr_dat[3] ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/res_mem_wr_dat[2] ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/res_mem_wr_dat[1] ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/res_mem_wr_dat[0] ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/res_mem_wr_addr[10] ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/res_mem_wr_addr[9] ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/res_mem_wr_addr[8] ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/res_mem_wr_addr[7] ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/res_mem_wr_addr[6] ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/res_mem_wr_addr[5] ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/res_mem_wr_addr[4] ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/res_mem_wr_addr[3] ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/res_mem_wr_addr[2] ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/res_mem_wr_addr[1] ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/res_mem_wr_addr[0] ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/res_mem_wr_pt[1] ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/res_mem_wr_pt[0] ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/resend_hp_act ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/tx_hdr_seq_num_dec[2] ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/tx_hdr_seq_num_dec[1] ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/tx_hdr_seq_num_dec[0] ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/resend_hp_num[4] ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/resend_hp_num[3] ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/resend_hp_num[2] ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/resend_hp_num[1] ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/resend_hp_num[0] ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/res_mem_rd_pt[1] ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/res_mem_rd_pt[0] ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/res_mem_rd_addr[10] ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/res_mem_rd_addr[9] ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/res_mem_rd_addr[8] ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/res_mem_rd_addr[7] ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/res_mem_rd_addr[6] ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/res_mem_rd_addr[5] ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/res_mem_rd_addr[4] ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/res_mem_rd_addr[3] ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/res_mem_rd_addr[2] ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/res_mem_rd_addr[1] ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/res_mem_rd_addr[0] ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/res_mem_rd_en ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/tx_res_req ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/tx_res_req_ack ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/res_mem_rd_dat[35] ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/res_mem_rd_dat[34] ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/res_mem_rd_dat[33] ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/res_mem_rd_dat[32] ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/res_mem_rd_dat[31] ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/res_mem_rd_dat[30] ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/res_mem_rd_dat[29] ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/res_mem_rd_dat[28] ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/res_mem_rd_dat[27] ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/res_mem_rd_dat[26] ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/res_mem_rd_dat[25] ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/res_mem_rd_dat[24] ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/res_mem_rd_dat[23] ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/res_mem_rd_dat[22] ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/res_mem_rd_dat[21] ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/res_mem_rd_dat[20] ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/res_mem_rd_dat[19] ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/res_mem_rd_dat[18] ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/res_mem_rd_dat[17] ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/res_mem_rd_dat[16] ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/res_mem_rd_dat[15] ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/res_mem_rd_dat[14] ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/res_mem_rd_dat[13] ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/res_mem_rd_dat[12] ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/res_mem_rd_dat[11] ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/res_mem_rd_dat[10] ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/res_mem_rd_dat[9] ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/res_mem_rd_dat[8] ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/res_mem_rd_dat[7] ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/res_mem_rd_dat[6] ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/res_mem_rd_dat[5] ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/res_mem_rd_dat[4] ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/res_mem_rd_dat[3] ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/res_mem_rd_dat[2] ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/res_mem_rd_dat[1] ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/res_mem_rd_dat[0] ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/res_mem_rd_dat_val ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/out_data_5[31] ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/out_data_5[30] ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/out_data_5[29] ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/out_data_5[28] ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/out_data_5[27] ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/out_data_5[26] ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/out_data_5[25] ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/out_data_5[24] ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/out_data_5[23] ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/out_data_5[22] ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/out_data_5[21] ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/out_data_5[20] ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/out_data_5[19] ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/out_data_5[18] ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/out_data_5[17] ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/out_data_5[16] ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/out_data_5[15] ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/out_data_5[14] ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/out_data_5[13] ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/out_data_5[12] ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/out_data_5[11] ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/out_data_5[10] ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/out_data_5[9] ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/out_data_5[8] ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/out_data_5[7] ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/out_data_5[6] ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/out_data_5[5] ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/out_data_5[4] ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/out_data_5[3] ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/out_data_5[2] ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/out_data_5[1] ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/out_data_5[0] ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/out_datak_5[3] ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/out_datak_5[2] ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/out_datak_5[1] ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/out_datak_5[0] ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/out_active_5 ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/tx_hdr_seq_num_dec_latch[2] ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/tx_hdr_seq_num_dec_latch[1] ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/tx_hdr_seq_num_dec_latch[0] ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/tx_lgood_empty ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/tx_lcrd_empty ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/send_hp_state[2] ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/send_hp_state[1] ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/send_hp_state[0] ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/send_lcmd_state[3] ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/send_lcmd_state[2] ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/send_lcmd_state[1] ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/send_lcmd_state[0] ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/tx_sel[2] ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/tx_sel[1] ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/tx_sel[0] ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/tx_lcrd_act ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/qc[7] ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/qc[6] ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/qc[5] ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/qc[4] ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/qc[3] ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/qc[2] ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/qc[1] ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/qc[0] ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/tx_lgood_act ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/res_state[2] ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/res_state[1] ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/res_state[0] ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/buf_out_dp_acked[2] ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/usb3_ep2_IN/buf_in_ready ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/usb3_ep2_IN/buf_in_commit ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/usb3_ep2_IN/buf_in_eob ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/usb3_ep2_IN/in_ep_rty ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/usb3_ep2_IN/buf_out_hasdata ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/usb3_ep2_IN/buf_out_eob ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/usb3_ep2_IN/buf_out_nump[4] ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/usb3_ep2_IN/buf_out_nump[3] ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/usb3_ep2_IN/buf_out_nump[2] ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/usb3_ep2_IN/buf_out_nump[1] ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/usb3_ep2_IN/buf_out_nump[0] ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/usb3_ep2_IN/buf_out_next_dp_ack_pt[3] ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/usb3_ep2_IN/buf_out_next_dp_ack_pt[2] ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/usb3_ep2_IN/buf_out_next_dp_ack_pt[1] ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/usb3_ep2_IN/buf_out_next_dp_ack_pt[0] ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/usb3_ep2_IN/buf_wt_ack_mem[15] ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/usb3_ep2_IN/buf_wt_ack_mem[14] ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/usb3_ep2_IN/buf_wt_ack_mem[13] ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/usb3_ep2_IN/buf_wt_ack_mem[12] ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/usb3_ep2_IN/buf_wt_ack_mem[11] ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/usb3_ep2_IN/buf_wt_ack_mem[10] ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/usb3_ep2_IN/buf_wt_ack_mem[9] ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/usb3_ep2_IN/buf_wt_ack_mem[8] ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/usb3_ep2_IN/buf_wt_ack_mem[7] ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/usb3_ep2_IN/buf_wt_ack_mem[6] ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/usb3_ep2_IN/buf_wt_ack_mem[5] ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/usb3_ep2_IN/buf_wt_ack_mem[4] ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/usb3_ep2_IN/buf_wt_ack_mem[3] ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/usb3_ep2_IN/buf_wt_ack_mem[2] ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/usb3_ep2_IN/buf_wt_ack_mem[1] ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/usb3_ep2_IN/buf_wt_ack_mem[0] ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/usb3_ep2_IN/buf_ready_mem[0] ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/usb3_ep2_IN/buf_ready_mem[1] ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/usb3_ep2_IN/buf_ready_mem[2] ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/usb3_ep2_IN/buf_ready_mem[3] ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/usb3_ep2_IN/buf_ready_mem[4] ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/usb3_ep2_IN/buf_ready_mem[5] ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/usb3_ep2_IN/buf_ready_mem[6] ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/usb3_ep2_IN/buf_ready_mem[7] ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/usb3_ep2_IN/buf_ready_mem[8] ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/usb3_ep2_IN/buf_ready_mem[9] ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/usb3_ep2_IN/buf_ready_mem[10] ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/usb3_ep2_IN/buf_ready_mem[11] ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/usb3_ep2_IN/buf_ready_mem[12] ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/usb3_ep2_IN/buf_ready_mem[13] ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/usb3_ep2_IN/buf_ready_mem[14] ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/usb3_ep2_IN/buf_ready_mem[15] ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/usb3_ep2_IN/buf_out_hasdata_mem[0] ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/usb3_ep2_IN/buf_out_hasdata_mem[1] ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/usb3_ep2_IN/buf_out_hasdata_mem[2] ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/usb3_ep2_IN/buf_out_hasdata_mem[3] ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/usb3_ep2_IN/buf_out_hasdata_mem[4] ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/usb3_ep2_IN/buf_out_hasdata_mem[5] ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/usb3_ep2_IN/buf_out_hasdata_mem[6] ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/usb3_ep2_IN/buf_out_hasdata_mem[7] ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/usb3_ep2_IN/buf_out_hasdata_mem[8] ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/usb3_ep2_IN/buf_out_hasdata_mem[9] ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/usb3_ep2_IN/buf_out_hasdata_mem[10] ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/usb3_ep2_IN/buf_out_hasdata_mem[11] ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/usb3_ep2_IN/buf_out_hasdata_mem[12] ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/usb3_ep2_IN/buf_out_hasdata_mem[13] ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/usb3_ep2_IN/buf_out_hasdata_mem[14] ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/usb3_ep2_IN/buf_out_hasdata_mem[15] ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/err_lbad_recv_latch ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/err_lbad_recv_latch_2 ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/usb3_ep2_IN/buf_out_pt[3] ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/usb3_ep2_IN/buf_out_pt[2] ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/usb3_ep2_IN/buf_out_pt[1] ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/usb3_ep2_IN/buf_out_pt[0] ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/usb3_ep2_IN/buf_in_pt[3] ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/usb3_ep2_IN/buf_in_pt[2] ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/usb3_ep2_IN/buf_in_pt[1] ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/usb3_ep2_IN/buf_in_pt[0] ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/usb3_ep2_IN/wt_ack_pt[3] ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/usb3_ep2_IN/wt_ack_pt[2] ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/usb3_ep2_IN/wt_ack_pt[1] ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3r/usb3_ep2_IN/wt_ack_pt[0] ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/tx_hp_act ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/err_hp_seq_latch ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/err_lgood_order_latch ,\USB30_Device_Controller_Top_inst/usb30_device_controller_inst/iu3l/tx_lgood_pop }),
    .clk_i(pclk)
);

endmodule
