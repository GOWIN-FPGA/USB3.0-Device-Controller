`define Q1_LN1
